��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�ű��k��'D��cd�w��i'OAWĎ(��./1b��w��д�nQ�(L	Ȉ���.0a��
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�{���_�<g��D+_�n��!�D-Fu����S�[��y: ��˘磋��w�����H���h=���D��F�omI	���������t���2�[�28�B�I:׷�F����"��/��\�vūx`��:�֡�\�<7�X�e�ʳ�A~�0 �i7�sp>7.~Ƨ����?2^�9�OI'�V�'n�^0o����y�]�$�R�n���=cv �ʆ�In��t��|׾&�@����[ƺTZ94���H��,k�w]��n0B��Fn^����7!�^ֻ��!� c�"�;���Y�lM�Ӻ��L�g�ֆ�F���\�vūx`��:�ވ�'��Ǵ�X�)Х��؊�K�H��\�v��wc�}�![ވ�'��Ǵϴ`�-2�ﻋ-�����S8�E�qVf>�A<t���j��Y�8%���Q�0�	�A�����<��z��}�����z���}��~�Q��eHmglS*��dO��(M�rUA3�v�~������]�!��Ȅ�I�� �/������!n}y���q���U�nPk���d`o����;v�~������]�!��	Ǹ�y85���*�t�<]���P�.�a(􆿳�����|�z�)�XGG�č�Y���S�)37J*u��l�M��ոi��<�g�T<�t�S��{l�f|�ό���.� *����h��|���kJ�!n}y���q���U�<��$R�08��������)��[6���9�dMbZ鎬�����%�M��>�h$G�����=����(�
t��Y�{'%s=ͱu��̦�"�K�b��Ub�ۙD^�V]��}R�wX��y�J�#z����ͩ^��8k>6s����]�!��	Ǹ�y85�������&H�[&-n�g��U-�eӥ+�V��b܉���i�kL�5N�6�vg;Je'���Xw��4L2�����c-(���X$�{�b�@IE�U��@�ڗe'��Q�$�yf��nͼ<�TD���9�,�w� �:&�sSs�Ǆo}|��XH�����,>$<�խ5�P�h=���D��F�omI	�������'�*3 �?��i_ U�`�w���2��@����跤="�3�j��'K���#<q!:�+0�|e|p�`��<����L�Y&��ѻ�p�$Y��C�tH'a�;,��R�BE�?7s�9���o��S8� j�(�3k��`y���pzl��a�I��Jt���[�L
�4x���e�+�rs�i�:�pdG��8p.������Y6�y!%O�T�\ ���|.�Tӏ��zw��;��,��c��d�٣��c�A�L'{Z�˗D�6���l ^�V]��}��ł�!r�dN�<@Iv���a_|���pzl��a�اQ��9M7s�9���o��S8��m�o�&i~G��;ؔa��-)��Cҷ��e�ˇ�h��]�Hlu���a'�<� \[	sqX��I�\�W�EC����F��Z鎬����Y�V��#q+~'%�ͫ 0�݊�,E��Tj� @>�Z鎬����Ԗ^Z�4q󕏜9���14�~�Xo.ݰB�u�9%�Z鎬�������(���O���EWI��X�)Х���[� Ag��g��U-�eɖ2��ن�'���ߌ[#(焋�Y�yv<�1������
�?<�yǯϷm���\��E��U���}h��R�Q��=f׿�������!N�2��_:��y$[|�h���X ��ʯÄ��@�����t��y�|�q���~�"����7Xa0~���;A���p�����|AW��ʗ&���MԲ������M�u�����;I4���i
E��l�1�ԀU%T3��W< slxSwP6h���X �=l�o �<�V|G/����Q*J�<I��%����$s�'fa�A�
��vޣ{b�'���V�,!2P510*���6�0)^�ګ�����p����nj��sR6�.�iGJ�����o5���jz��j�(�2I�Sr����a!��h����0>��r��kGQ��l�4��H���0�0�h��#g�k�����x^6���[�L
ú�@�Z�\�����p�!a�bS펓$�R�n���M�a(􆿳��J���J6j�"Hs�U��Y���G��:!���v�H�~����Iu���r�pΚ�w]�L�� �0���E�+a�G3�u]˴�����x_��s�֙���C��f5�%��)f��20�	�>�� �~A�s�|����3-T}�p~G��;ؔa��-)��Cҷ��e[�� <7S�*���X�#Gw6�E��0Tm56���l ^�V]��}R�wX�Ձc������,!���[��2���2R=@�R�BE�?q��g�kD�w43��"�,�&�L4⭦Ϛ|�.qh;��|B�g��rB��y{�הr6�T��B_C�Z������=���>|�(�O��u����+P�W�躩�[��ɶ0h�5e���{t�XE�j$���X��WG ���j�!�	?:��E�Q�%]n9��Mv!���x�%�`�ʾ�Oߤy6��}@!;��Va�ir��dc�@�E��g@�M��.�X�y����.Oe���"X}�a&�s$- ��/"��и�]+z�@_-�H���J�1���۪	�}a4������J�>�_C�Z���&Q�[���Q�6D��x�Ӷ	F�ukc��f)�%\��s�o.;��f:_�A�M6'	|�+��?�d���&��v�<����@DO]�5����V�m�������։EF�6���l �4�9ܡ��#g�k��g?	��o�y����Rb�ɵ�Zr��s�{�����d����5��P,�%[Z럡~�H�B� ��~���4M̍���Qw�c4~Nrg�d�h��`�ѧ$u�{�6��5�ź�q9+t�}�G=X���8�P��Gh�1 :�[�d��-��!���0I52z���a��M�"w�wP��d�p�,�����n�Ak����
�u��٫fL����x{^4��*m-}ʙLY�>QR��Q��#�K4�d��rLF��ٹ�F���$�R�n���Mڰ���k�l׏�����MFi��|��wØ�ߤ\Dvk��u�R8H�[���R'cf���:ڢ�[��p.������Y6�y!%O?�d���&��G=X��cx������g~�/��>�Y`�}^AH?�d���&�n<�y{�הr.}e�'�K�5~2Qr�B�M�5�Y����+>Q ����)c�4��>.g�K:+>�+5�X��������Ut�\����=5Z'pǘ���Mv!���x�\�G�����Qf=��1���`��@w���H��j�Ï��	p8,3s"X��WG ���D�$0�	���SQ����:|-M�O��~�΢�u�L���7����̡L��)�I>|�(�O��l�;V��p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�φ��<�6��9�8;eM���w����E� ����՝��z|�6��1�I�I���мC%��2�S�OߙYĸ-r9p��-��o�>���mB�GOu"��c������,!��b��8!
��z%�ژ�(|k��|���X�7QZ����x#� P!���.�_�8��$�R�n���Mڂf>x�:	�E�&�y++���Ã8�4��Q>��\d:0�g��MY����̎,������)�PuS��_��<Q�G�`f���s}��$Ck;�a�<d��[&�$*�9U<���Hn
V~$�c��Z�q(�a�df;[�����a�z6��\d:0�g���D8�I�/xR��\&4��Ȝx��y���-M�O��~Ӿ9�d�L��di���̋'Q�|����\��~U��-�R5���,"~������[��x��y�o���9V�S^NLH�&7G֨˜��Cи�]+z�@��jO�(cc�}���Fo|k�LbJ�1���K���L���߸��S�Ȍ���Y���_� 
��,������=<�6>'r {�Q�%��)f��'T���'�&�8C�����8Χ�
��Uq��1��XNLH�&7�NjX�U�6j�"Hs�}����V:\�2*ޢƍgR��r��ܦ_����{���28E)CO���&�L4⭦��n�z�t?�d���&�n<�y{�הr.}e�'�K�5~2QrǷ�:h�(n�.�p������?��9)����M��k$��"T N��r*�D�$0�Qw�c4~Nrg�d��%�z�J��	���SQ���嫋�T���Hp9��m��;�����6�h,�@#o�]�ʄ�m�Թ���pY)�/����l*8��dUt�\�͋�߬JoNLH�&7������mo���SK�%_C�Z���5��s�kχ�n|,�Rn
V~$@�	��K��/B結�JA�d��rLF��ٹ�F���^���EqJ�1��씑�:��KY׏�����M����!2�͞nOY� �U�O��Dx�A�A=���g��K���|_b9 ��%��)f��'T���'��O�Jc�H_C�Z����܊����ZD�[?���ѧ$u�{�6��5�źm���?�e�yyg��yY|�6��1�I�I���мC%��2�SRu�y��C��hhjq�>.�)����:�'�V��	��yte�wqs*��7�E�Um1�H���W�w��fD��`}�8�`�ҧ��?�d���&��:�=�R�0�1�]  #��P	�qB�o!f�	�Ĳ��Bf���{^��6G����f�iC��{Q[��n���yXEƈ�o!f�	�Ĳ��Bf���rs�(�̴Y�{'%s�ui�铊���͚�2�TZ94���}Ņ��<��DΦ��t�x�=����H��efm�0z�cUL���ޤ�Y5�`]�n�p�V|����26���l ŃP�|�A6(�u<*~G��;ؔ��Νd[�*�������h�6Q�7���yoZ�P/Ȗa�N�����E� ���$�R�n���M�au'�;�iݘ��C_�矻�vt2��EyS�쇥�_��o�s(㷾���E.t�