module psw (
    input clk, g, g_en,
    output reg gf
);

// gf��ʼֵΪ0
initial begin
    gf = 1'b0;
end

// ��ʱ���½��ظ��¼Ĵ���
always @(negedge clk) begin
    if (g_en)
        gf <= g; // ��� g_en Ϊ 1�����Ĵ�����ֵ����Ϊ�����ź� g
end

endmodule
