��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5�h��%��Xcbp��'����Q4KҲ��r�D� �m�'�t�חEʭ�3�Jld��q�G�~��Z2��˝1~OT������oPY̅���c�PƐt
׫�J��q{�f��a�:&�>��s�z+/�c�Z�J
_䆼�\�v�����{�{\J�yG����y��\�vť���ҧ`�S�*H������=t����w���@�|��].��'���Xwd�n]Nِ����_H;a(􆿳���A�b,�my$�N���Uە��GV��y�&_3#ڸZ鎬����D�OBp�b}��BB϶q��{l�f|�ό���.Ӳ�[O�"���Ig`i�ҋX����@�ڗe'��E4�Mʸ|��].��'���Xw�-X��-���Ig`i�ҋX����@�ڗe'�@.�>�ȼ�|��].��'���Xw����UA����Ig`i7G#+���[H�����2��~��o�b�x�'�6LE�EYZ/���)֨9 >�j��O0E>�������fHa��!A{�H]�%�Iߎn?�e"�2ao
r��FE���r#�9l$���޸�����C�O"I��MjX��k���`���F(ĕL2	X�vb�)�S�����]�c.��'1����1\���k�e1i��Q,�&d���ݚev3Y�IkT˱ ��O�������]�U�����8�o��@�<�qؚ��L�NG�>)�����7������7�� �����R=�;@R��Ω�dBj#/����@$˺/tw�ԝD=��٭@�FϟQ�-i�`�g``FD�e3>�ƙ�Ǘ���mC��XH�����wI�d��`���1�E��)֨9 E3����=E�EYZ/�@�L0�6#����"'W�9�p��y��9��L����Lo�I��'��恭�h�I��'�%�e���Ĕ^ֻ��X�x%}�����
D�5tm�c�oL�~j�F},M�5����`K�����svfY������;5B5Y+���o�(�)��;U��tm�c�oL�������FTVP��b�M:�8U(�d�٣��c�A�L'��y�!�;&����˚�T�\ �����j�|�z#:rQ��q�X�G[��;ۂ���cY�~�"���ʷ��1�(ʌ�N�M8�U����t��h~��J����^Mf���9���q���U�pzl��a��i��؂ۃ�y�wjאﻋ-�����S8�l��`�_gi�.�!����Wy����`y����s��d�\��MN����!I/�������A��X�@�5��6�l��sХ+�:R 8*!Ē\��c�PƐt
�20)�_�5�e��a)�m�d�so�}a�C�ub;�;���A���g?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��Le��	I���]�HЦ��EMW!���4m~�����c-�z��~��D:ǯ3�4���X�E��	�'�J���U�2Gޣסe� <���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+�S�AZL�0hs�A_	�K�o[��mU;լ^<���X�E��j I�ƹ�+��nV]J�l�!y�Y�RZ/�+"�����}q�����>��9����W��l����4�n���xǊ��i�������}���7��./�>.���k1O#�+T���t_-Z��T�\ ���s��r-���CE�ow�2@���z�������v齅�"Dh\�n):��Bo�A;h�F$�Μ��VK)q7p�5jG�P�֯�=k�Rm���}d�����s��B��Kj%��A5'��|��V�4v!4���ts2����,J!�w:��������Ut�\�A��R�ߋQ"���_޾I�_�*@Z������/dN�<@Iv��nt=:�-���)z�$8Fs�<���Hn
V~$E��>����^(�<<���Hn
V~$E$Ԣ���[m�(��k8���i�|.N,�z_M?ą����ȳ��(���5zCo�����.��24��i��Q�J���8��Z��������d�*�e�qb"q|��˓#�����t�)�A�ސ���d�w#��\�ސ���'d��i�)J�1��쌳���������"O��tm�c�oL�;U�Qb���|�B��6Yd2��΃����~���vX��N��24��L���Y�nȗ;Øh�ه� �4�<+�����UrD�zU�����f���NRP`��!;��I#��p�-a�D͢�����.�B�R���>_�ryO#��!�Y��N������%��T�\ ��Ǫ�v�/P)�6�=�#��11�g��U-�eMg.6�kcw���n���k��i�}0.���s�5�e��0UJ�1����ݾ-/�uu��ڿ׏�����M��ܐ�}�&��������}���:!�׿M?S{V*(��N�ߎ���#-!N�'�y�G