-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.


LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY TRIBUF_a8237 IS
    PORT (
        in1 : IN std_logic;
        oe  : IN std_logic;
        y   : OUT std_logic);
END TRIBUF_a8237;

ARCHITECTURE behavior OF TRIBUF_a8237 IS
BEGIN
    PROCESS (in1, oe)
    BEGIN
        IF oe'EVENT THEN
            IF oe = '0' THEN
                y <= TRANSPORT 'Z'  ;
            ELSIF oe = '1' THEN
                y <= TRANSPORT in1  ;
            END IF;
        ELSIF oe = '1' THEN
            y <= TRANSPORT in1  ;
        END IF;
    END PROCESS;
END behavior;

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DFF_a8237 IS
    PORT (
      	 d   : IN std_logic;
      	 clk : IN std_logic;
      	 clrn: IN std_logic;
      	 prn : IN std_logic;
      	 q   : OUT std_logic := '0');
END DFF_a8237;

ARCHITECTURE behavior OF DFF_a8237 IS
BEGIN

    PROCESS (clk, clrn, prn)
        VARIABLE result : std_logic := '0';
    BEGIN
        ASSERT NOT (prn = '0' AND clrn = '0')
            REPORT " prn and clrn both '0' on DFF"
            SEVERITY Warning;

        IF prn = '0' AND clrn = '1' THEN
            result := '1';
        ELSIF prn = '1' AND clrn = '0' THEN
            result := '0';
        ELSIF rising_edge(clk) THEN
            IF d = '1' OR d = '0' THEN
                result := d;
            END IF;
        END IF;

        IF result /= 'X' THEN
            q <= TRANSPORT result  ;
        END IF;

    END PROCESS;
END behavior;

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY FILTER_a8237 IS
    PORT (
        in1 : IN std_logic;
        y: OUT std_logic);
END FILTER_a8237;

ARCHITECTURE behavior OF FILTER_a8237 IS
BEGIN

    y <= in1;
END behavior;

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE work.tribuf_a8237;
USE work.dff_a8237;
USE work.filter_a8237;

ENTITY a8237 IS
    PORT (
      ain : IN std_logic_vector(3 downto 0);
      dbin : IN std_logic_vector(7 downto 0);
      dreq : IN std_logic_vector(3 downto 0);
      aout : OUT std_logic_vector(7 downto 0);
      dack : OUT std_logic_vector(3 downto 0);
      dbout : OUT std_logic_vector(7 downto 0);
      clk : IN std_logic;
      hlda : IN std_logic;
      ncs : IN std_logic;
      neopin : IN std_logic;
      niorin : IN std_logic;
      niowin : IN std_logic;
      ready : IN std_logic;
      reset : IN std_logic;
      adstb : OUT std_logic;
      aen : OUT std_logic;
      dben : OUT std_logic;
      dmaenable : OUT std_logic;
      hrq : OUT std_logic;
      neopout : OUT std_logic;
      niorout : OUT std_logic;
      niowout : OUT std_logic;
      nmemr : OUT std_logic;
      nmemw : OUT std_logic);
END a8237;

ARCHITECTURE Version_1_0 OF a8237 IS

SIGNAL gnd : std_logic := '0';
SIGNAL vcc : std_logic := '1';
SIGNAL
    n_153, n_154, n_155, n_156, n_157, a_G956, n_159, n_160, n_161, n_162,
          n_163, n_164, a_G1027, n_166, n_167, n_168, n_169, n_170, n_171,
          a_G200, n_173, n_174, n_175, n_176, n_177, n_178, a_G186, n_180,
          n_181, n_182, n_183, n_184, n_185, a_G993, n_187, n_188, n_189,
          n_190, n_191, n_192, a_G917, n_194, n_195, n_196, n_197, n_198,
          n_199, a_G142, n_201, n_202, n_203, n_204, n_205, n_206, a_G1389,
          n_208, n_209, n_210, n_211, n_212, n_213, a_G503, n_215, n_216,
          n_217, n_218, n_219, n_220, a_G502, n_222, n_223, n_224, n_225,
          n_226, n_227, a_G1464, n_229, n_230, n_231, n_232, n_233, n_234,
          a_G1463, n_236, n_237, n_238, n_239, n_240, n_241, a_LC7_D18, n_243,
          n_244, n_245, n_246, n_247, n_248, a_LC7_C17, n_250, n_251, n_252,
          n_253, n_254, n_255, a_LC4_C16, n_257, n_258, n_259, n_260, n_261,
          n_262, a_LC2_C24, n_264, n_265, n_266, n_267, n_268, n_269, a_LC1_C16,
          n_271, n_272, n_273, n_274, n_275, n_276, a_LC3_F6, n_278, n_279,
          n_280, n_281, n_282, n_283, a_LC4_F10, n_285, n_286, n_287, n_288,
          n_289, n_290, a_LC5_D27, n_292, n_293, n_294, n_295, n_296, n_297,
          a_SNMEMW, n_299, n_300, n_301, n_302, n_303, n_304, a_SNMEMR_aNOT,
          n_306, n_307, n_308, n_309, n_310, n_311, a_SNIOWOUT, n_313, n_314,
          n_315, n_316, n_317, n_318, a_SNIOROUT, n_320, n_321, n_322, n_323,
          n_324, n_325, a_SNEOPOUT_aNOT, n_327, n_328, n_329, n_330, n_331,
          n_332, a_SHRQ, n_334, n_335, n_336, n_337, n_338, n_339, a_SAEN_aNOT,
          n_341, n_342, n_343, n_344, n_345, n_346, a_SDBEN, n_348, n_349,
          n_350, n_351, n_352, n_353, a_LC6_B16_aNOT, n_355, n_356, n_357,
          n_358, n_359, n_360, a_SADSTB, n_362, a_SCH2BWORDOUT_F3_G, a_SCH2BWORDOUT_F3_G_aCLRN,
          a_EQ1030, n_371, n_372, n_373, a_N2574_aNOT, n_375, n_377, n_378,
          n_379, n_380, n_381, a_SCH2BWORDOUT_F3_G_aCLK, a_SCH0BWORDOUT_F4_G,
          a_SCH0BWORDOUT_F4_G_aCLRN, a_EQ903, n_391, n_392, n_393, a_N2578_aNOT,
          n_395, n_397, n_398, n_399, n_400, n_401, a_SCH0BWORDOUT_F4_G_aCLK,
          a_SCH3BWORDOUT_F4_G, a_SCH3BWORDOUT_F4_G_aCLRN, a_EQ1095, n_410,
          n_411, n_412, a_N2572_aNOT, n_414, n_415, n_416, n_417, n_418, n_419,
          a_SCH3BWORDOUT_F4_G_aCLK, a_SCH2BWORDOUT_F4_G, a_SCH2BWORDOUT_F4_G_aCLRN,
          a_EQ1031, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435,
          n_436, a_SCH2BWORDOUT_F4_G_aCLK, a_SCH1BWORDOUT_F4_G, a_SCH1BWORDOUT_F4_G_aCLRN,
          a_EQ967, n_445, n_446, n_447, a_N2576_aNOT, n_449, n_450, n_451,
          n_452, n_453, n_454, a_SCH1BWORDOUT_F4_G_aCLK, a_N2352, a_EQ556,
          n_458, n_459, n_460, n_462, n_463, n_465, n_466, n_468, n_469, n_471,
          a_N2585_aNOT, a_EQ638, n_474, n_475, n_476, n_477, n_478, a_LC3_D22,
          n_480, a_SCH1BAROUT_F12_G, a_SCH1BAROUT_F12_G_aCLRN, a_EQ959, n_488,
          n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, a_SCH1BAROUT_F12_G_aCLK,
          a_SCH1BAROUT_F13_G, a_SCH1BAROUT_F13_G_aCLRN, a_EQ960, n_505, n_506,
          n_507, n_508, n_510, n_511, n_512, n_513, n_514, a_SCH1BAROUT_F13_G_aCLK,
          a_SCH2BWORDOUT_F6_G, a_SCH2BWORDOUT_F6_G_aCLRN, a_EQ1033, n_523,
          n_524, n_525, n_526, n_528, n_529, n_530, n_531, n_532, a_SCH2BWORDOUT_F6_G_aCLK,
          a_SCH1BWORDOUT_F6_G, a_SCH1BWORDOUT_F6_G_aCLRN, a_EQ969, n_541,
          n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, a_SCH1BWORDOUT_F6_G_aCLK,
          a_SCH0BWORDOUT_F6_G, a_SCH0BWORDOUT_F6_G_aCLRN, a_EQ905, n_558,
          n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, a_SCH0BWORDOUT_F6_G_aCLK,
          a_N77_aNOT, a_EQ194, n_570, n_571, n_572, n_573, n_574, n_575, n_576,
          n_577, n_578, n_579, a_N2583_aNOT, a_EQ636, n_582, n_583, n_584,
          n_585, n_586, n_587, a_SCH2BAROUT_F14_G, a_SCH2BAROUT_F14_G_aCLRN,
          a_EQ1025, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602,
          n_603, a_SCH2BAROUT_F14_G_aCLK, a_SCH1BAROUT_F14_G, a_SCH1BAROUT_F14_G_aCLRN,
          a_EQ961, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619,
          n_620, a_SCH1BAROUT_F14_G_aCLK, a_SCH1BWORDOUT_F7_G, a_SCH1BWORDOUT_F7_G_aCLRN,
          a_EQ970, n_629, n_630, n_631, n_632, n_634, n_635, n_636, n_637,
          n_638, a_SCH1BWORDOUT_F7_G_aCLK, a_N2573_aNOT, a_EQ626, n_642, n_643,
          n_644, bytepointer, n_646, n_647, a_N87, n_649, n_650, a_N2347,
          n_652, a_SCH3BWORDOUT_F11_G, a_SCH3BWORDOUT_F11_G_aCLRN, a_EQ1102,
          n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, a_SCH3BWORDOUT_F11_G_aCLK,
          a_SCH1BWORDOUT_F11_G, a_SCH1BWORDOUT_F11_G_aCLRN, a_EQ974, n_677,
          n_678, n_679, a_N2577_aNOT, n_681, n_682, n_683, n_684, n_685, n_686,
          a_SCH1BWORDOUT_F11_G_aCLK, a_SCH2BWORDOUT_F11_G, a_SCH2BWORDOUT_F11_G_aCLRN,
          a_EQ1038, n_695, n_696, n_697, n_698, a_N62_aNOT, n_700, n_701,
          n_702, n_703, n_704, n_705, n_706, n_707, n_708, a_SCH2BWORDOUT_F11_G_aCLK,
          a_SCH0BWORDOUT_F11_G, a_SCH0BWORDOUT_F11_G_aCLRN, a_EQ910, n_717,
          n_718, n_719, n_720, a_N2353, n_722, n_723, n_724, n_725, n_726,
          n_727, n_728, n_729, n_730, a_SCH0BWORDOUT_F11_G_aCLK, a_SCH3BWORDOUT_F12_G,
          a_SCH3BWORDOUT_F12_G_aCLRN, a_EQ1103, n_739, n_740, n_741, n_742,
          n_743, n_744, n_745, n_746, n_747, a_SCH3BWORDOUT_F12_G_aCLK, a_SCH0BWORDOUT_F12_G,
          a_SCH0BWORDOUT_F12_G_aCLRN, a_EQ911, n_756, n_757, n_758, n_759,
          n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, a_SCH0BWORDOUT_F12_G_aCLK,
          a_SCH2BWORDOUT_F12_G, a_SCH2BWORDOUT_F12_G_aCLRN, a_EQ1039, n_777,
          n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787,
          n_788, n_789, a_SCH2BWORDOUT_F12_G_aCLK, a_SCH1BWORDOUT_F12_G, a_SCH1BWORDOUT_F12_G_aCLRN,
          a_EQ975, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805,
          n_806, a_SCH1BWORDOUT_F12_G_aCLK, a_SCH3BWORDOUT_F2_G, a_SCH3BWORDOUT_F2_G_aCLRN,
          a_EQ1093, n_815, n_816, n_817, n_818, n_820, n_821, n_822, n_823,
          n_824, a_SCH3BWORDOUT_F2_G_aCLK, a_SCH2BWORDOUT_F2_G, a_SCH2BWORDOUT_F2_G_aCLRN,
          a_EQ1029, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840,
          n_841, a_SCH2BWORDOUT_F2_G_aCLK, a_SCH3BWORDOUT_F14_G, a_SCH3BWORDOUT_F14_G_aCLRN,
          a_EQ1105, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857,
          n_858, a_SCH3BWORDOUT_F14_G_aCLK, a_SCH1BWORDOUT_F14_G, a_SCH1BWORDOUT_F14_G_aCLRN,
          a_EQ977, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874,
          n_875, a_SCH1BWORDOUT_F14_G_aCLK, a_SCH2BWORDOUT_F14_G, a_SCH2BWORDOUT_F14_G_aCLRN,
          a_EQ1041, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891,
          n_892, n_893, n_894, n_895, n_896, a_SCH2BWORDOUT_F14_G_aCLK, a_SCH0BWORDOUT_F14_G,
          a_SCH0BWORDOUT_F14_G_aCLRN, a_EQ913, n_905, n_906, n_907, n_908,
          n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, a_SCH0BWORDOUT_F14_G_aCLK,
          a_LC1_C22, a_EQ024, n_921, n_922, n_923, a_N3554, n_925, a_N3556,
          n_927, n_928, n_929, a_N3555, n_931, n_932, n_933, n_934, n_935,
          a_LC4_A3, a_EQ192, n_938, n_939, n_940, n_941, n_942, n_943, n_944,
          n_945, a_N2563_aNOT, a_EQ616, n_948, n_949, n_950, n_951, n_952,
          n_953, n_954, n_955, a_N70, a_N70_aIN, n_958, n_959, n_960, a_N820,
          n_962, a_N822, n_964, a_N821, n_966, a_N823, n_968, a_N71_aNOT,
          a_EQ190, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978,
          n_979, n_980, a_LC1_B23_aNOT, a_EQ574, n_983, n_984, n_985, n_986,
          n_987, n_988, n_989, n_990, a_N2361, a_EQ562, n_993, n_994, n_995,
          n_996, n_997, n_998, a_N1584, a_EQ472, n_1001, n_1002, n_1003, n_1004,
          n_1005, n_1006, n_1007, n_1008, a_N2557, a_N2557_aIN, n_1011, n_1012,
          n_1013, n_1014, n_1015, a_N1164_aNOT, a_EQ374, n_1018, n_1019, n_1020,
          n_1021, n_1022, n_1023, n_1024, n_1025, a_N2598_aNOT, a_EQ647, n_1028,
          n_1029, n_1030, a_SCHANNEL_F1_G, n_1032, n_1033, a_SCHANNEL_F0_G,
          n_1035, a_N2591, a_N2591_aIN, n_1038, n_1039, n_1040, n_1041, a_SCOMMANDREG_F0_G,
          n_1043, a_N2531, a_N2531_aIN, n_1046, n_1047, n_1048, n_1049, n_1050,
          a_N2374, a_EQ568, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058,
          n_1059, n_1060, n_1061, n_1062, a_N2408_aNOT, a_EQ579, n_1065, n_1066,
          n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074,
          n_1075, n_1076, n_1077, n_1078, a_N68_aNOT, a_EQ188, n_1081, n_1082,
          n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090,
          a_LC4_B25_aNOT, a_LC4_B25_aNOT_aIN, n_1093, n_1094, n_1095, n_1096,
          n_1097, a_N67_aNOT, a_EQ187, n_1100, n_1101, n_1102, n_1103, n_1104,
          n_1105, n_1106, n_1107, n_1108, n_1109, a_N2356, a_EQ559, n_1112,
          n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120,
          n_1121, a_N1592, a_N1592_aIN, n_1124, n_1125, n_1126, n_1127, n_1128,
          n_1129, a_N1566, a_EQ465, n_1132, n_1133, n_1134, n_1135, n_1136,
          n_1137, n_1138, n_1139, a_N2358, a_EQ560, n_1142, n_1143, n_1144,
          n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, a_LC8_B20,
          a_EQ476, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160,
          n_1161, n_1162, n_1163, n_1164, a_N1588, a_N1588_aIN, n_1167, n_1168,
          n_1169, n_1170, n_1171, n_1172, a_N88_aNOT, a_EQ197, n_1175, n_1176,
          n_1177, n_1178, n_1179, n_1180, a_N2377, a_EQ570, n_1183, n_1184,
          n_1185, n_1186, n_1187, n_1188, a_LC4_E22, a_EQ580, n_1191, n_1192,
          n_1193, n_1194, a_SCH1MODEREG_F1_G, n_1196, n_1197, n_1198, a_SCH3MODEREG_F1_G,
          n_1200, a_N2376, a_EQ569, n_1203, n_1204, n_1205, n_1206, n_1207,
          n_1208, a_LC6_E22, a_EQ582, n_1211, n_1212, n_1213, a_SCH2MODEREG_F0_G,
          n_1215, a_SCH1MODEREG_F0_G, n_1217, n_1218, n_1219, n_1220, n_1221,
          n_1222, n_1223, n_1224, n_1225, n_1226, a_LC5_E22, a_EQ583, n_1229,
          n_1230, n_1231, a_SCH0MODEREG_F0_G, n_1233, a_SCH3MODEREG_F0_G,
          n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242,
          n_1243, n_1244, a_LC6_E10, a_EQ581, n_1247, n_1248, n_1249, n_1250,
          a_SCH0MODEREG_F1_G, n_1252, n_1253, n_1254, a_SCH2MODEREG_F1_G,
          n_1256, a_N1589, a_EQ478, n_1259, n_1260, n_1261, n_1262, n_1263,
          n_1264, n_1265, n_1266, n_1267, n_1268, a_N1580_aNOT, a_EQ468, n_1271,
          n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279,
          n_1280, a_SNMEMR_aNOT_aIN, n_1282, n_1283, n_1284, n_1285, n_1286,
          n_1287, a_N1180, a_EQ385, n_1290, n_1291, n_1292, n_1293, a_SCH1WRDCNTREG_F2_G,
          n_1295, n_1296, n_1297, a_SCH0WRDCNTREG_F2_G, n_1299, a_LC4_C6,
          a_EQ386, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308,
          n_1309, a_LC2_C6, a_EQ384, n_1312, n_1313, n_1314, n_1315, a_SCH2WRDCNTREG_F2_G,
          n_1317, n_1318, n_1319, a_SCH3WRDCNTREG_F2_G, n_1321, a_LC1_C6,
          a_EQ383, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330,
          n_1331, a_N3554_aCLRN, a_EQ850, n_1338, n_1339, n_1340, n_1341,
          startdma, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349,
          n_1350, a_N3554_aCLK, a_LC7_C22, a_EQ023, n_1354, n_1355, n_1356,
          n_1357, n_1358, n_1359, n_1360, n_1361, a_LC4_C27, a_EQ361, n_1364,
          n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372,
          a_LC6_C27, a_EQ363, n_1375, n_1376, n_1377, n_1378, a_SCH1WRDCNTREG_F1_G,
          n_1380, n_1381, n_1382, a_SCH3WRDCNTREG_F1_G, n_1384, a_LC2_C27,
          a_EQ364, n_1387, n_1388, n_1389, n_1390, a_SCH2WRDCNTREG_F1_G, n_1392,
          n_1393, n_1394, a_SCH0WRDCNTREG_F1_G, n_1396, a_N1139, a_EQ365,
          n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406,
          a_LC5_C27, a_EQ362, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414,
          n_1415, n_1416, n_1417, n_1418, a_N3555_aCLRN, a_EQ851, n_1425,
          n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433,
          n_1434, n_1435, n_1436, a_N3555_aCLK, a_LC1_C21, a_EQ025, n_1440,
          n_1441, n_1442, n_1443, a_N3553, n_1445, n_1446, n_1447, n_1448,
          n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456,
          a_LC7_C15, a_EQ253, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464,
          n_1465, n_1466, a_LC5_C15, a_EQ254, n_1469, n_1470, n_1471, n_1472,
          a_SCH1WRDCNTREG_F3_G, n_1474, n_1475, n_1476, a_SCH0WRDCNTREG_F3_G,
          n_1478, a_N491_aNOT, a_EQ255, n_1481, n_1482, n_1483, n_1484, n_1485,
          n_1486, n_1487, n_1488, a_LC5_C14, a_EQ257, n_1491, n_1492, n_1493,
          n_1494, a_SCH3WRDCNTREG_F3_G, n_1496, n_1497, n_1498, a_SCH2WRDCNTREG_F3_G,
          n_1500, a_LC1_C15, a_EQ256, n_1503, n_1504, n_1505, n_1506, n_1507,
          n_1508, n_1509, n_1510, a_N3553_aCLRN, a_EQ849, n_1517, n_1518,
          n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526,
          n_1527, n_1528, a_N3553_aCLK, a_SCH2BAROUT_F8_G, a_SCH2BAROUT_F8_G_aCLRN,
          a_EQ1019, n_1537, n_1538, n_1539, n_1540, n_1542, n_1543, n_1544,
          n_1545, n_1546, a_SCH2BAROUT_F8_G_aCLK, a_SCH3BWORDOUT_F8_G, a_SCH3BWORDOUT_F8_G_aCLRN,
          a_EQ1099, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561,
          n_1562, n_1563, a_SCH3BWORDOUT_F8_G_aCLK, a_N2354_aNOT, a_N2354_aNOT_aIN,
          n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, a_N2586,
          a_N2586_aIN, n_1576, n_1577, n_1578, a_LC6_D6, n_1580, n_1581, a_N2587_aNOT,
          a_EQ640, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, a_SCH0BAROUT_F8_G,
          a_SCH0BAROUT_F8_G_aCLRN, a_EQ891, n_1597, n_1598, n_1599, n_1600,
          n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608,
          n_1609, a_SCH0BAROUT_F8_G_aCLK, a_N2348, a_EQ554, n_1613, n_1614,
          n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622,
          a_N2581_aNOT, a_EQ632, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630,
          a_SCH3BAROUT_F8_G, a_SCH3BAROUT_F8_G_aCLRN, a_EQ1083, n_1638, n_1639,
          n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, a_SCH3BAROUT_F8_G_aCLK,
          a_SCH0BWORDOUT_F8_G, a_SCH0BWORDOUT_F8_G_aCLRN, a_EQ907, n_1655,
          n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663,
          n_1664, n_1665, n_1666, n_1667, a_SCH0BWORDOUT_F8_G_aCLK, a_SCH1BAROUT_F8_G,
          a_SCH1BAROUT_F8_G_aCLRN, a_EQ955, n_1676, n_1677, n_1678, n_1679,
          n_1680, n_1681, n_1682, n_1683, n_1684, a_SCH1BAROUT_F8_G_aCLK,
          a_SCH2BWORDOUT_F8_G, a_SCH2BWORDOUT_F8_G_aCLRN, a_EQ1035, n_1693,
          n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701,
          n_1702, n_1703, n_1704, n_1705, a_SCH2BWORDOUT_F8_G_aCLK, a_SCH1BWORDOUT_F8_G,
          a_SCH1BWORDOUT_F8_G_aCLRN, a_EQ971, n_1714, n_1715, n_1716, n_1717,
          n_1718, n_1719, n_1720, n_1721, n_1722, a_SCH1BWORDOUT_F8_G_aCLK,
          a_SCH3BWORDOUT_F0_G, a_SCH3BWORDOUT_F0_G_aCLRN, a_EQ1091, n_1731,
          n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739,
          a_SCH3BWORDOUT_F0_G_aCLK, a_SCH0BWORDOUT_F0_G, a_SCH0BWORDOUT_F0_G_aCLRN,
          a_EQ899, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754,
          n_1755, n_1756, a_SCH0BWORDOUT_F0_G_aCLK, a_SCH2BWORDOUT_F0_G, a_SCH2BWORDOUT_F0_G_aCLRN,
          a_EQ1027, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771,
          n_1772, n_1773, a_SCH2BWORDOUT_F0_G_aCLK, a_LC8_D12, a_EQ516, n_1777,
          n_1778, n_1779, n_1780, a_SCH0WRDCNTREG_F0_G, n_1782, n_1783, n_1784,
          a_SCH1WRDCNTREG_F0_G, n_1786, a_N1867_aNOT, a_EQ515, n_1789, n_1790,
          n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798,
          n_1799, n_1800, n_1801, a_LC5_D12, a_EQ514, n_1804, n_1805, n_1806,
          n_1807, a_SCH3WRDCNTREG_F0_G, n_1809, n_1810, n_1811, n_1812, a_LC6_D12,
          a_EQ513, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821,
          a_SCH2WRDCNTREG_F0_G, n_1823, a_N3556_aCLRN, a_EQ852, n_1830, n_1831,
          n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839,
          n_1840, n_1841, a_N3556_aCLK, a_SCH3BAROUT_F9_G, a_SCH3BAROUT_F9_G_aCLRN,
          a_EQ1084, n_1850, n_1851, n_1852, n_1853, n_1855, n_1856, n_1857,
          n_1858, n_1859, a_SCH3BAROUT_F9_G_aCLK, a_SCH2BAROUT_F9_G, a_SCH2BAROUT_F9_G_aCLRN,
          a_EQ1020, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874,
          n_1875, n_1876, a_SCH2BAROUT_F9_G_aCLK, a_SCH0BAROUT_F9_G, a_SCH0BAROUT_F9_G_aCLRN,
          a_EQ892, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891,
          n_1892, n_1893, a_SCH0BAROUT_F9_G_aCLK, a_LC3_C13, a_EQ036, n_1897,
          n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905,
          n_1906, a_LC8_F13_aNOT, a_LC8_F13_aNOT_aIN, n_1909, n_1910, n_1911,
          n_1912, a_N3552, n_1914, a_N3551, n_1916, a_N3550, n_1918, a_LC4_A13_aNOT,
          a_LC4_A13_aNOT_aIN, n_1921, n_1922, n_1923, n_1924, a_N3549, n_1926,
          a_N3548, n_1928, a_N3547, n_1930, a_LC1_A20_aNOT, a_LC1_A20_aNOT_aIN,
          n_1933, n_1934, n_1935, n_1936, a_N3546, n_1938, a_N3545, n_1940,
          a_N3544, n_1942, a_LC3_E16_aNOT, a_LC3_E16_aNOT_aIN, n_1945, n_1946,
          n_1947, n_1948, a_N3543, n_1950, a_N3542, n_1952, a_N2539, a_N2539_aIN,
          n_1955, n_1956, n_1957, n_1958, a_N3541, n_1960, a_LC1_B12, a_EQ1164,
          n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970,
          n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978,
          n_1979, n_1980, a_EQ1163, n_1982, n_1983, n_1984, n_1985, n_1986,
          n_1987, n_1988, n_1989, n_1990, n_1991, a_N57_aNOT, a_EQ181, n_1994,
          n_1995, n_1996, n_1997, n_1998, n_1999, a_N825, n_2001, a_N2528,
          a_N2528_aIN, n_2004, n_2005, n_2006, n_2007, a_SCH3MODEREG_F2_G,
          n_2009, a_N965, a_EQ331, n_2012, n_2013, n_2014, n_2015, n_2016,
          n_2017, a_N1095, a_N1095_aIN, n_2020, n_2021, n_2022, n_2023, n_2024,
          a_LC3_C4, a_EQ832, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032,
          n_2033, n_2034, n_2035, n_2036, a_N1046_aNOT, a_N1046_aNOT_aIN,
          n_2039, n_2040, n_2041, a_SCH3BWORDOUT_F1_G, n_2043, n_2044, a_N1094,
          a_N1094_aIN, n_2047, n_2048, n_2049, n_2050, n_2051, a_SCH3WRDCNTREG_F1_G_aCLRN,
          a_EQ1114, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064,
          n_2065, n_2066, n_2067, a_SCH3WRDCNTREG_F1_G_aCLK, a_N2558_aNOT,
          a_EQ613, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077,
          n_2078, n_2079, a_LC1_C12, a_EQ771, n_2082, n_2083, n_2084, n_2085,
          n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093,
          a_LC2_C12, a_EQ772, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101,
          n_2102, n_2103, a_N2525, a_N2525_aIN, n_2106, n_2107, n_2108, n_2109,
          a_SCH0MODEREG_F2_G, n_2111, a_SCH0WRDCNTREG_F1_G_aCLRN, a_EQ922,
          n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, a_SCH0BWORDOUT_F1_G,
          n_2125, n_2126, n_2127, a_SCH0WRDCNTREG_F1_G_aCLK, a_N2559_aNOT,
          a_EQ614, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137,
          n_2138, n_2139, n_2140, a_N2526, a_N2526_aIN, n_2143, n_2144, n_2145,
          n_2146, a_SCH1MODEREG_F2_G, n_2148, a_N2595, a_N2595_aIN, n_2151,
          n_2152, n_2153, n_2154, n_2155, a_LC7_D26, a_LC7_D26_aIN, n_2158,
          n_2159, n_2160, n_2161, n_2162, a_LC6_A25, a_EQ793, n_2165, n_2166,
          n_2167, n_2168, n_2169, n_2170, a_SCH1BWORDOUT_F1_G, n_2172, n_2173,
          a_N433, a_N433_aIN, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181,
          n_2182, a_N460, a_N460_aIN, n_2185, n_2186, n_2187, n_2188, n_2189,
          a_SCH1WRDCNTREG_F1_G_aCLRN, a_EQ986, n_2196, n_2197, n_2198, n_2199,
          n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, a_SCH1WRDCNTREG_F1_G_aCLK,
          a_N2560_aNOT, a_EQ615, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214,
          a_N2527, a_N2527_aIN, n_2217, n_2218, n_2219, n_2220, a_SCH2MODEREG_F2_G,
          n_2222, a_N756, a_N756_aIN, n_2225, n_2226, n_2227, n_2228, n_2229,
          a_LC2_C18, a_EQ812, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237,
          n_2238, n_2239, n_2240, n_2241, a_N797, a_N797_aIN, n_2244, n_2245,
          n_2246, a_SCH2BWORDOUT_F1_G, n_2248, n_2249, a_N858, a_N858_aIN,
          n_2252, n_2253, n_2254, n_2255, n_2256, a_SCH2WRDCNTREG_F1_G_aCLRN,
          a_EQ1050, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269,
          n_2270, n_2271, n_2272, a_SCH2WRDCNTREG_F1_G_aCLK, a_LC1_A13, a_EQ028,
          n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283,
          n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291,
          a_LC3_A7, a_EQ758, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299,
          n_2300, n_2301, a_SCH0WRDCNTREG_F9_G, n_2303, n_2304, n_2305, n_2306,
          a_LC4_A7, a_EQ759, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314,
          n_2315, n_2316, a_SCH0WRDCNTREG_F9_G_aCLRN, a_EQ930, n_2323, n_2324,
          n_2325, n_2326, n_2327, n_2328, a_SCH0BWORDOUT_F9_G, n_2330, n_2331,
          n_2332, a_SCH0WRDCNTREG_F9_G_aCLK, a_LC2_E12, a_LC2_E12_aIN, n_2336,
          n_2337, n_2338, n_2339, n_2340, a_LC3_A25, a_EQ782, n_2343, n_2344,
          n_2345, n_2346, a_SCH1WRDCNTREG_F9_G, n_2348, n_2349, a_SCH1BWORDOUT_F9_G,
          n_2351, n_2352, a_N636_aNOT, a_N636_aNOT_aIN, n_2355, n_2356, n_2357,
          n_2358, n_2359, n_2360, n_2361, a_SCH1WRDCNTREG_F9_G_aCLRN, a_EQ994,
          n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375,
          n_2376, n_2377, a_SCH1WRDCNTREG_F9_G_aCLK, a_LC1_A7, a_EQ803, n_2381,
          n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, a_SCH2WRDCNTREG_F9_G,
          n_2390, n_2391, n_2392, n_2393, a_LC2_A7, a_EQ804, n_2396, n_2397,
          n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, a_SCH2WRDCNTREG_F9_G_aCLRN,
          a_EQ1058, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, a_SCH2BWORDOUT_F9_G,
          n_2417, n_2418, n_2419, a_SCH2WRDCNTREG_F9_G_aCLK, a_SCH1BAROUT_F9_G,
          a_SCH1BAROUT_F9_G_aCLRN, a_EQ956, n_2428, n_2429, n_2430, n_2431,
          n_2432, n_2433, n_2434, n_2435, n_2436, a_SCH1BAROUT_F9_G_aCLK,
          a_SCH3BWORDOUT_F9_G, a_SCH3BWORDOUT_F9_G_aCLRN, a_EQ1100, n_2445,
          n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453,
          a_SCH3BWORDOUT_F9_G_aCLK, a_SCH0BWORDOUT_F2_G, a_SCH0BWORDOUT_F2_G_aCLRN,
          a_EQ901, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468,
          n_2469, n_2470, a_SCH0BWORDOUT_F2_G_aCLK, a_SCH2BAROUT_F10_G, a_SCH2BAROUT_F10_G_aCLRN,
          a_EQ1021, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485,
          n_2486, n_2487, a_SCH2BAROUT_F10_G_aCLK, a_SCH3BWORDOUT_F10_G, a_SCH3BWORDOUT_F10_G_aCLRN,
          a_EQ1101, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502,
          n_2503, n_2504, a_SCH3BWORDOUT_F10_G_aCLK, a_SCH3BAROUT_F10_G, a_SCH3BAROUT_F10_G_aCLRN,
          a_EQ1085, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519,
          n_2520, n_2521, a_SCH3BAROUT_F10_G_aCLK, a_SCH2BWORDOUT_F10_G, a_SCH2BWORDOUT_F10_G_aCLRN,
          a_EQ1037, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536,
          n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, a_SCH2BWORDOUT_F10_G_aCLK,
          a_SCH1BAROUT_F10_G, a_SCH1BAROUT_F10_G_aCLRN, a_EQ957, n_2551, n_2552,
          n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, a_SCH1BAROUT_F10_G_aCLK,
          a_SCH0BWORDOUT_F10_G, a_SCH0BWORDOUT_F10_G_aCLRN, a_EQ909, n_2568,
          n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576,
          n_2577, n_2578, n_2579, n_2580, a_SCH0BWORDOUT_F10_G_aCLK, a_SCH0BAROUT_F10_G,
          a_SCH0BAROUT_F10_G_aCLRN, a_EQ893, n_2589, n_2590, n_2591, n_2592,
          n_2593, n_2594, n_2595, n_2596, n_2597, a_SCH0BAROUT_F10_G_aCLK,
          a_SCH2BAROUT_F11_G, a_SCH2BAROUT_F11_G_aCLRN, a_EQ1022, n_2606,
          n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614,
          a_SCH2BAROUT_F11_G_aCLK, a_SCH3BAROUT_F11_G, a_SCH3BAROUT_F11_G_aCLRN,
          a_EQ1086, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629,
          n_2630, n_2631, a_SCH3BAROUT_F11_G_aCLK, a_SCH0BAROUT_F11_G, a_SCH0BAROUT_F11_G_aCLRN,
          a_EQ894, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646,
          n_2647, n_2648, a_SCH0BAROUT_F11_G_aCLK, a_SCH1BAROUT_F11_G, a_SCH1BAROUT_F11_G_aCLRN,
          a_EQ958, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663,
          n_2664, n_2665, a_SCH1BAROUT_F11_G_aCLK, a_LC1_C10, a_EQ767, n_2669,
          n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, a_LC3_C10,
          a_EQ768, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685,
          n_2686, a_SCH0WRDCNTREG_F3_G_aCLRN, a_EQ924, n_2693, n_2694, n_2695,
          n_2696, n_2697, n_2698, a_SCH0BWORDOUT_F3_G, n_2700, n_2701, n_2702,
          a_SCH0WRDCNTREG_F3_G_aCLK, a_LC2_C22, a_EQ790, n_2706, n_2707, n_2708,
          n_2709, n_2710, n_2711, n_2712, n_2713, a_LC5_C22, a_EQ791, n_2716,
          n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, a_SCH1WRDCNTREG_F3_G_aCLRN,
          a_EQ988, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, a_SCH1BWORDOUT_F3_G,
          n_2737, n_2738, n_2739, a_SCH1WRDCNTREG_F3_G_aCLK, a_LC2_C7, a_EQ810,
          n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750,
          n_2751, n_2752, a_N808, a_N808_aIN, n_2755, n_2756, n_2757, n_2758,
          n_2759, a_SCH2WRDCNTREG_F3_G_aCLRN, a_EQ1052, n_2766, n_2767, n_2768,
          n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, a_SCH2WRDCNTREG_F3_G_aCLK,
          a_SCH3BWORDOUT_F3_G, a_SCH3BWORDOUT_F3_G_aCLRN, a_EQ1094, n_2784,
          n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792,
          a_SCH3BWORDOUT_F3_G_aCLK, a_LC1_C3, a_EQ765, n_2796, n_2797, n_2798,
          n_2799, n_2800, n_2801, n_2802, a_SCH0WRDCNTREG_F4_G, n_2804, a_LC2_C3,
          a_EQ766, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813,
          n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, a_SCH0WRDCNTREG_F4_G_aCLRN,
          a_EQ925, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832,
          n_2833, n_2834, a_SCH0WRDCNTREG_F4_G_aCLK, a_LC2_C1, a_EQ829, n_2838,
          n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846,
          a_SCH3WRDCNTREG_F4_G, n_2848, a_N1037_aNOT, a_EQ344, n_2851, n_2852,
          n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860,
          a_SCH3WRDCNTREG_F4_G_aCLRN, a_EQ1117, n_2867, n_2868, n_2869, n_2870,
          n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, a_SCH3WRDCNTREG_F4_G_aCLK,
          a_LC4_C18, a_EQ809, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885,
          n_2886, n_2887, n_2888, a_SCH2WRDCNTREG_F4_G, n_2890, a_N815, a_EQ304,
          n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900,
          n_2901, n_2902, a_SCH2WRDCNTREG_F4_G_aCLRN, a_EQ1053, n_2909, n_2910,
          n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918,
          a_SCH2WRDCNTREG_F4_G_aCLK, a_LC5_F4, a_EQ788, n_2922, n_2923, n_2924,
          n_2925, n_2926, n_2927, n_2928, a_SCH1WRDCNTREG_F4_G, n_2930, a_LC6_F4,
          a_EQ789, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939,
          n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, a_SCH1WRDCNTREG_F4_G_aCLRN,
          a_EQ989, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958,
          n_2959, n_2960, a_SCH1WRDCNTREG_F4_G_aCLK, a_SCH2BAROUT_F12_G, a_SCH2BAROUT_F12_G_aCLRN,
          a_EQ1023, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975,
          n_2976, n_2977, a_SCH2BAROUT_F12_G_aCLK, a_SCH0BAROUT_F12_G, a_SCH0BAROUT_F12_G_aCLRN,
          a_EQ895, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992,
          n_2993, n_2994, a_SCH0BAROUT_F12_G_aCLK, a_SCH3BAROUT_F12_G, a_SCH3BAROUT_F12_G_aCLRN,
          a_EQ1087, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009,
          n_3010, n_3011, a_SCH3BAROUT_F12_G_aCLK, a_SCH0BWORDOUT_F5_G, a_SCH0BWORDOUT_F5_G_aCLRN,
          a_EQ904, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026,
          n_3027, n_3028, a_SCH0BWORDOUT_F5_G_aCLK, a_SCH3BWORDOUT_F5_G, a_SCH3BWORDOUT_F5_G_aCLRN,
          a_EQ1096, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043,
          n_3044, n_3045, a_SCH3BWORDOUT_F5_G_aCLK, a_SCH1BWORDOUT_F5_G, a_SCH1BWORDOUT_F5_G_aCLRN,
          a_EQ968, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060,
          n_3061, n_3062, a_SCH1BWORDOUT_F5_G_aCLK, a_SCH2BWORDOUT_F5_G, a_SCH2BWORDOUT_F5_G_aCLRN,
          a_EQ1032, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077,
          n_3078, n_3079, a_SCH2BWORDOUT_F5_G_aCLK, a_SCH0BWORDOUT_F13_G,
          a_SCH0BWORDOUT_F13_G_aCLRN, a_EQ912, n_3088, n_3089, n_3090, n_3091,
          n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099,
          n_3100, a_SCH0BWORDOUT_F13_G_aCLK, a_SCH3BWORDOUT_F13_G, a_SCH3BWORDOUT_F13_G_aCLRN,
          a_EQ1104, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115,
          n_3116, n_3117, a_SCH3BWORDOUT_F13_G_aCLK, a_SCH1BWORDOUT_F13_G,
          a_SCH1BWORDOUT_F13_G_aCLRN, a_EQ976, n_3126, n_3127, n_3128, n_3129,
          n_3130, n_3131, n_3132, n_3133, n_3134, a_SCH1BWORDOUT_F13_G_aCLK,
          a_SCH2BWORDOUT_F13_G, a_SCH2BWORDOUT_F13_G_aCLRN, a_EQ1040, n_3143,
          n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151,
          n_3152, n_3153, n_3154, n_3155, a_SCH2BWORDOUT_F13_G_aCLK, a_SCH2BAROUT_F13_G,
          a_SCH2BAROUT_F13_G_aCLRN, a_EQ1024, n_3164, n_3165, n_3166, n_3167,
          n_3168, n_3169, n_3170, n_3171, n_3172, a_SCH2BAROUT_F13_G_aCLK,
          a_SCH0BAROUT_F13_G, a_SCH0BAROUT_F13_G_aCLRN, a_EQ896, n_3181, n_3182,
          n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, a_SCH0BAROUT_F13_G_aCLK,
          a_SCH3BAROUT_F13_G, a_SCH3BAROUT_F13_G_aCLRN, a_EQ1088, n_3198,
          n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206,
          a_SCH3BAROUT_F13_G_aCLK, a_LC7_F24, a_EQ807, n_3210, n_3211, n_3212,
          n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, a_SCH2WRDCNTREG_F6_G,
          n_3220, a_LC7_F13, a_EQ026, n_3223, n_3224, n_3225, n_3226, n_3227,
          n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235,
          n_3236, n_3237, n_3238, a_N832_aNOT, a_N832_aNOT_aIN, n_3241, n_3242,
          n_3243, n_3244, n_3245, n_3246, a_SCH2WRDCNTREG_F6_G_aCLRN, a_EQ1055,
          n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260,
          n_3261, n_3262, a_SCH2WRDCNTREG_F6_G_aCLK, a_LC5_F27, a_EQ827, n_3266,
          n_3267, n_3268, n_3269, n_3270, n_3271, a_SCH3BWORDOUT_F6_G, n_3273,
          n_3274, a_N1066, a_EQ349, n_3277, n_3278, n_3279, n_3280, n_3281,
          n_3282, n_3283, a_SCH3WRDCNTREG_F6_G, n_3285, a_SCH3WRDCNTREG_F6_G_aCLRN,
          a_EQ1119, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298,
          n_3299, a_SCH3WRDCNTREG_F6_G_aCLK, a_LC1_F4, a_EQ785, n_3303, n_3304,
          n_3305, n_3306, n_3307, n_3308, n_3309, a_SCH1WRDCNTREG_F6_G, n_3311,
          a_LC2_F4, a_EQ786, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319,
          n_3320, n_3321, a_SCH1WRDCNTREG_F6_G_aCLRN, a_EQ991, n_3328, n_3329,
          n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, a_SCH1WRDCNTREG_F6_G_aCLK,
          a_LC2_F8, a_EQ762, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345,
          n_3346, a_SCH0WRDCNTREG_F6_G, n_3348, a_LC4_F8, a_EQ763, n_3351,
          n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, a_SCH0WRDCNTREG_F6_G_aCLRN,
          a_EQ927, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371,
          n_3372, n_3373, a_SCH0WRDCNTREG_F6_G_aCLK, a_SCH0BAROUT_F14_G, a_SCH0BAROUT_F14_G_aCLRN,
          a_EQ897, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388,
          n_3389, n_3390, a_SCH0BAROUT_F14_G_aCLK, a_SCH3BAROUT_F14_G, a_SCH3BAROUT_F14_G_aCLRN,
          a_EQ1089, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405,
          n_3406, n_3407, a_SCH3BAROUT_F14_G_aCLK, a_SCH3BWORDOUT_F7_G, a_SCH3BWORDOUT_F7_G_aCLRN,
          a_EQ1098, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422,
          n_3423, n_3424, a_SCH3BWORDOUT_F7_G_aCLK, a_SCH2BWORDOUT_F7_G, a_SCH2BWORDOUT_F7_G_aCLRN,
          a_EQ1034, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439,
          n_3440, n_3441, a_SCH2BWORDOUT_F7_G_aCLK, a_SCH0BWORDOUT_F7_G, a_SCH0BWORDOUT_F7_G_aCLRN,
          a_EQ906, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456,
          n_3457, n_3458, a_SCH0BWORDOUT_F7_G_aCLK, a_SCH2BAROUT_F15_G, a_SCH2BAROUT_F15_G_aCLRN,
          a_EQ1026, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473,
          n_3474, n_3475, a_SCH2BAROUT_F15_G_aCLK, a_SCH0BAROUT_F15_G, a_SCH0BAROUT_F15_G_aCLRN,
          a_EQ898, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490,
          n_3491, n_3492, a_SCH0BAROUT_F15_G_aCLK, a_SCH3BAROUT_F15_G, a_SCH3BAROUT_F15_G_aCLRN,
          a_EQ1090, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507,
          n_3508, n_3509, a_SCH3BAROUT_F15_G_aCLK, a_SCH1BAROUT_F15_G, a_SCH1BAROUT_F15_G_aCLRN,
          a_EQ962, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524,
          n_3525, n_3526, a_SCH1BAROUT_F15_G_aCLK, a_LC5_A20, a_EQ029, n_3530,
          n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538,
          n_3539, n_3540, n_3541, a_LC4_A22, a_EQ820, n_3544, n_3545, n_3546,
          n_3547, n_3548, n_3549, n_3550, a_SH3WRDCNTREG_F11_G, n_3552, a_LC3_A22,
          a_EQ821, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561,
          n_3562, a_SH3WRDCNTREG_F11_G_aCLRN, a_EQ1152, n_3569, n_3570, n_3571,
          n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, a_SH3WRDCNTREG_F11_G_aCLK,
          a_LC5_A11, a_EQ778, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586,
          n_3587, a_SH1WRDCNTREG_F11_G, n_3589, a_LC3_A11, a_EQ779, n_3592,
          n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, a_SH1WRDCNTREG_F11_G_aCLRN,
          a_EQ1140, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612,
          n_3613, n_3614, a_SH1WRDCNTREG_F11_G_aCLK, a_LC4_F26, a_EQ799, n_3618,
          n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, a_SH2WRDCNTREG_F11_G,
          n_3627, n_3628, n_3629, n_3630, a_LC5_F26, a_EQ800, n_3633, n_3634,
          n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, a_SH2WRDCNTREG_F11_G_aCLRN,
          a_EQ1146, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653,
          n_3654, n_3655, a_SH2WRDCNTREG_F11_G_aCLK, a_LC5_A22, a_EQ756, n_3659,
          n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, a_SH0WRDCNTREG_F11_G,
          n_3668, n_3669, n_3670, n_3671, a_LC6_A22, a_EQ757, n_3674, n_3675,
          n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, a_SH0WRDCNTREG_F11_G_aCLRN,
          a_EQ1134, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694,
          n_3695, n_3696, a_SH0WRDCNTREG_F11_G_aCLK, a_LC6_A20, a_EQ030, n_3700,
          n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708,
          n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, a_LC3_A21,
          a_EQ818, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724,
          a_SH3WRDCNTREG_F12_G, n_3726, a_LC4_A21, a_EQ819, n_3729, n_3730,
          n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, a_SH3WRDCNTREG_F12_G_aCLRN,
          a_EQ1153, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749,
          n_3750, n_3751, a_SH3WRDCNTREG_F12_G_aCLK, a_LC1_A8, a_EQ754, n_3755,
          n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, a_SH0WRDCNTREG_F12_G,
          n_3764, n_3765, n_3766, n_3767, a_LC2_A8, a_EQ755, n_3770, n_3771,
          n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, a_SH0WRDCNTREG_F12_G_aCLRN,
          a_EQ1135, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790,
          n_3791, n_3792, a_SH0WRDCNTREG_F12_G_aCLK, a_LC3_A14, a_EQ797, n_3796,
          n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, a_SH2WRDCNTREG_F12_G,
          n_3805, n_3806, n_3807, n_3808, a_LC2_A14, a_EQ798, n_3811, n_3812,
          n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, a_SH2WRDCNTREG_F12_G_aCLRN,
          a_EQ1147, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831,
          n_3832, n_3833, a_SH2WRDCNTREG_F12_G_aCLK, a_LC1_A11, a_EQ776, n_3837,
          n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, a_SH1WRDCNTREG_F12_G,
          n_3845, a_LC2_A11, a_EQ777, n_3848, n_3849, n_3850, n_3851, n_3852,
          n_3853, n_3854, n_3855, a_SH1WRDCNTREG_F12_G_aCLRN, a_EQ1141, n_3862,
          n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870,
          a_SH1WRDCNTREG_F12_G_aCLK, a_SCH0BWORDOUT_F15_G, a_SCH0BWORDOUT_F15_G_aCLRN,
          a_EQ914, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885,
          n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, a_SCH0BWORDOUT_F15_G_aCLK,
          a_SCH1BWORDOUT_F15_G, a_SCH1BWORDOUT_F15_G_aCLRN, a_EQ978, n_3900,
          n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908,
          a_SCH1BWORDOUT_F15_G_aCLK, a_SCH2BWORDOUT_F15_G, a_SCH2BWORDOUT_F15_G_aCLRN,
          a_EQ1042, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923,
          n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, a_SCH2BWORDOUT_F15_G_aCLK,
          a_SCH3BWORDOUT_F15_G, a_SCH3BWORDOUT_F15_G_aCLRN, a_EQ1106, n_3938,
          n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946,
          a_SCH3BWORDOUT_F15_G_aCLK, a_LC6_E16, a_EQ031, n_3950, n_3951, n_3952,
          n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960,
          n_3961, a_LC6_E5, a_EQ352, n_3964, n_3965, n_3966, n_3967, n_3968,
          n_3969, n_3970, a_SH3WRDCNTREG_F14_G, n_3972, a_LC5_E5, a_EQ646,
          n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982,
          a_SH3WRDCNTREG_F14_G_aCLRN, a_EQ1155, n_3989, n_3990, n_3991, n_3992,
          n_3993, n_3994, n_3995, n_3996, n_3997, a_SH3WRDCNTREG_F14_G_aCLK,
          a_N869_aNOT, a_EQ318, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006,
          n_4007, a_SH1WRDCNTREG_F14_G, n_4009, a_LC7_E19, a_EQ316, n_4012,
          n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, a_SH1WRDCNTREG_F14_G_aCLRN,
          a_EQ1143, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032,
          n_4033, n_4034, a_SH1WRDCNTREG_F14_G_aCLK, a_LC8_E4, a_EQ314, n_4038,
          n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, a_SH2WRDCNTREG_F14_G,
          n_4047, n_4048, n_4049, n_4050, a_LC7_E4, a_EQ323, n_4053, n_4054,
          n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, a_SH2WRDCNTREG_F14_G_aCLRN,
          a_EQ1149, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073,
          n_4074, n_4075, a_SH2WRDCNTREG_F14_G_aCLK, a_LC2_E13, a_EQ750, n_4079,
          n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, a_SH0WRDCNTREG_F14_G,
          n_4088, n_4089, n_4090, n_4091, a_LC3_E13, a_EQ751, n_4094, n_4095,
          n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, a_SH0WRDCNTREG_F14_G_aCLRN,
          a_EQ1137, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114,
          n_4115, n_4116, a_SH0WRDCNTREG_F14_G_aCLK, a_LC2_C25, a_EQ399, n_4120,
          n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, a_N1296_aNOT,
          a_EQ409, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136,
          n_4137, n_4138, n_4139, n_4140, n_4141, a_N1280, a_EQ398, n_4144,
          n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, a_N1279,
          a_EQ397, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160,
          n_4161, n_4162, n_4163, a_LC3_C25, a_EQ400, n_4166, n_4167, n_4168,
          n_4169, n_4170, n_4171, n_4172, n_4173, a_N3552_aCLRN, a_EQ848,
          n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, n_4187,
          n_4188, n_4189, n_4190, n_4191, a_N3552_aCLK, a_LC6_F16, a_EQ268,
          n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202,
          n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210,
          a_LC4_F16, a_EQ267, n_4213, n_4214, n_4215, n_4216, a_SCH1WRDCNTREG_F5_G,
          n_4218, n_4219, n_4220, a_SCH0WRDCNTREG_F5_G, n_4222, a_N522_aNOT,
          a_EQ264, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231,
          n_4232, a_LC3_F16, a_EQ266, n_4235, n_4236, n_4237, n_4238, a_SCH2WRDCNTREG_F5_G,
          n_4240, n_4241, n_4242, n_4243, a_LC1_F16, a_EQ265, n_4246, n_4247,
          n_4248, n_4249, n_4250, n_4251, n_4252, a_SCH3WRDCNTREG_F5_G, n_4254,
          a_N3551_aCLRN, a_EQ847, n_4261, n_4262, n_4263, n_4264, n_4265,
          n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, a_N3551_aCLK,
          a_LC6_F13, a_EQ505, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281,
          n_4282, n_4283, a_LC5_F13, a_EQ504, n_4286, n_4287, n_4288, n_4289,
          n_4290, n_4291, n_4292, n_4293, a_N1764_aNOT, a_EQ506, n_4296, n_4297,
          n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, a_LC1_F13, a_EQ503,
          n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313,
          a_LC2_F13, a_EQ502, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321,
          n_4322, n_4323, a_N3550_aCLRN, a_EQ846, n_4330, n_4331, n_4332,
          n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340,
          n_4341, a_N3550_aCLK, a_LC1_E11, a_EQ518, n_4345, n_4346, n_4347,
          n_4348, a_SCH0MODEREG_F3_G, n_4350, n_4351, n_4352, a_SCH1MODEREG_F3_G,
          n_4354, a_N1879_aNOT, a_EQ517, n_4357, n_4358, n_4359, n_4360, n_4361,
          n_4362, n_4363, n_4364, n_4365, n_4366, a_LC1_E1, a_EQ589, n_4369,
          n_4370, n_4371, n_4372, a_SCH3MODEREG_F3_G, n_4374, n_4375, n_4376,
          a_SCH2MODEREG_F3_G, n_4378, a_N2529, a_EQ590, n_4381, n_4382, n_4383,
          n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, a_N2530_aNOT,
          a_EQ591, n_4393, n_4394, n_4395, a_SCOMMANDREG_F1_G, n_4397, n_4398,
          n_4399, a_N757, a_N757_aIN, n_4402, n_4403, n_4404, n_4405, n_4406,
          a_LC2_C14, a_EQ002, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414,
          n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422,
          n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430,
          n_4431, n_4432, n_4433, n_4434, a_LC6_C14, a_LC6_C14_aIN, n_4437,
          n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445,
          n_4446, n_4447, a_LC3_C14, a_EQ019, n_4450, n_4451, n_4452, n_4453,
          n_4454, n_4455, n_4456, n_4457, a_LC4_C14, a_EQ021, n_4460, n_4461,
          n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469,
          n_4470, n_4471, n_4472, n_4473, n_4474, a_LC7_C14, a_EQ020, n_4477,
          n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485,
          n_4486, n_4487, n_4488, n_4489, a_LC1_F26, a_EQ003, n_4492, n_4493,
          n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501,
          n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509,
          n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517,
          a_LC4_F20, a_LC4_F20_aIN, n_4520, n_4521, n_4522, n_4523, n_4524,
          n_4525, n_4526, n_4527, n_4528, n_4529, n_4530, a_LC6_F20, a_EQ017,
          n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540,
          a_LC6_F15, a_EQ016, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548,
          n_4549, n_4550, n_4551, n_4552, n_4553, a_LC4_F15, a_EQ004, n_4556,
          n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, a_LC1_F15,
          a_EQ015, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572,
          n_4573, a_LC2_F14, a_EQ295, n_4576, n_4577, n_4578, n_4579, n_4580,
          n_4581, a_SADDRESSOUT_F8_G, n_4583, n_4584, n_4585, n_4586, n_4587,
          n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595,
          n_4596, n_4597, n_4598, a_LC1_F14, a_EQ713, n_4601, n_4602, n_4603,
          n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, a_SCH2ADDRREG_F8_G,
          n_4611, a_SCH2ADDRREG_F8_G_aCLRN, a_EQ1003, n_4618, n_4619, n_4620,
          n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628,
          n_4629, a_SCH2ADDRREG_F8_G_aCLK, a_LC5_D1, a_EQ223, n_4633, n_4634,
          n_4635, n_4636, n_4637, n_4638, n_4639, a_SCH3WRDCNTREG_F8_G, n_4641,
          a_LC6_D17, a_EQ027, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649,
          n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, a_LC6_D1, a_EQ224,
          n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665,
          a_SCH3WRDCNTREG_F8_G_aCLRN, a_EQ1121, n_4672, n_4673, n_4674, n_4675,
          n_4676, n_4677, n_4678, n_4679, n_4680, a_SCH3WRDCNTREG_F8_G_aCLK,
          a_N2548, a_EQ605, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689,
          n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697,
          n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705,
          n_4706, a_LC1_F7, a_EQ659, n_4709, n_4710, n_4711, n_4712, n_4713,
          n_4714, n_4715, a_SCH0ADDRREG_F8_G, n_4717, a_LC2_F7, a_EQ660, n_4720,
          n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, a_SCH0ADDRREG_F8_G_aCLRN,
          a_EQ875, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740,
          n_4741, n_4742, a_SCH0ADDRREG_F8_G_aCLK, a_LC5_F12, a_EQ330, n_4746,
          n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754,
          n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, n_4762,
          n_4763, n_4764, n_4765, n_4766, n_4767, a_LC2_F12, a_EQ738, n_4770,
          n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778,
          a_SCH3ADDRREG_F8_G, n_4780, a_SCH3ADDRREG_F8_G_aCLRN, a_EQ1067,
          n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794,
          n_4795, n_4796, n_4797, n_4798, a_SCH3ADDRREG_F8_G_aCLK, a_LC6_D10,
          a_EQ432, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808,
          n_4809, a_SCH0WRDCNTREG_F8_G, n_4811, n_4812, n_4813, n_4814, a_LC8_D10,
          a_EQ433, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823,
          n_4824, a_SCH0WRDCNTREG_F8_G_aCLRN, a_EQ929, n_4831, n_4832, n_4833,
          n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, a_SCH0WRDCNTREG_F8_G_aCLK,
          a_N1553, a_N1553_aIN, n_4843, n_4844, n_4845, n_4846, n_4847, a_LC7_F18,
          a_EQ460, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856,
          n_4857, n_4858, a_SCH1ADDRREG_F8_G, n_4860, a_SCH1ADDRREG_F8_G_aCLRN,
          a_EQ939, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873,
          n_4874, n_4875, n_4876, n_4877, n_4878, a_SCH1ADDRREG_F8_G_aCLK,
          a_N689_aNOT, a_EQ284, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887,
          n_4888, n_4889, a_SCH2WRDCNTREG_F8_G, n_4891, n_4892, n_4893, n_4894,
          a_LC3_D7, a_EQ805, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902,
          n_4903, n_4904, a_SCH2WRDCNTREG_F8_G_aCLRN, a_EQ1057, n_4911, n_4912,
          n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, a_SCH2WRDCNTREG_F8_G_aCLK,
          a_N357_aNOT, a_EQ236, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928,
          n_4929, a_SCH1WRDCNTREG_F8_G, n_4931, a_LC3_D1, a_EQ783, n_4934,
          n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, a_SCH1WRDCNTREG_F8_G_aCLRN,
          a_EQ993, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954,
          n_4955, n_4956, a_SCH1WRDCNTREG_F8_G_aCLK, a_LC3_D2, a_EQ833, n_4960,
          n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968,
          n_4969, a_N1033_aNOT, a_N1033_aNOT_aIN, n_4972, n_4973, n_4974,
          n_4975, n_4976, a_SCH3WRDCNTREG_F0_G_aCLRN, a_EQ1113, n_4983, n_4984,
          n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992,
          a_SCH3WRDCNTREG_F0_G_aCLK, a_N241_aNOT, a_EQ220, n_4996, n_4997,
          n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, a_LC2_D16, a_EQ773,
          n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013,
          a_SCH0WRDCNTREG_F0_G_aCLRN, a_EQ921, n_5020, n_5021, n_5022, n_5023,
          n_5024, n_5025, n_5026, n_5027, n_5028, a_SCH0WRDCNTREG_F0_G_aCLK,
          a_LC4_D20, a_EQ813, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037,
          n_5038, n_5039, n_5040, n_5041, a_N805, a_N805_aIN, n_5044, n_5045,
          n_5046, n_5047, n_5048, a_SCH2WRDCNTREG_F0_G_aCLRN, a_EQ1049, n_5055,
          n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063,
          n_5064, a_SCH2WRDCNTREG_F0_G_aCLK, a_LC7_D16, a_EQ794, n_5068, n_5069,
          n_5070, n_5071, n_5072, n_5073, a_SCH1BWORDOUT_F0_G, n_5075, n_5076,
          a_N435, a_N435_aIN, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084,
          a_SCH1WRDCNTREG_F0_G_aCLRN, a_EQ985, n_5091, n_5092, n_5093, n_5094,
          n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, a_SCH1WRDCNTREG_F0_G_aCLK,
          a_LC1_F10, a_EQ014, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109,
          n_5110, n_5111, n_5112, n_5113, n_5114, a_LC3_A2, a_EQ005, n_5117,
          n_5118, n_5119, n_5120, a_SADDRESSOUT_F9_G, n_5122, n_5123, n_5124,
          n_5125, a_LC4_A15, a_EQ736, n_5128, n_5129, n_5130, n_5131, n_5132,
          n_5133, n_5134, n_5135, a_SCH3ADDRREG_F9_G, n_5137, n_5138, n_5139,
          n_5140, a_LC6_A15, a_EQ737, n_5143, n_5144, n_5145, n_5146, n_5147,
          n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155,
          a_SCH3ADDRREG_F9_G_aCLRN, a_EQ1068, n_5162, n_5163, n_5164, n_5165,
          n_5166, n_5167, n_5168, n_5169, n_5170, a_SCH3ADDRREG_F9_G_aCLK,
          a_LC4_A16, a_EQ711, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179,
          n_5180, a_SCH2ADDRREG_F9_G, n_5182, a_LC6_A16, a_EQ712, n_5185,
          n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193,
          n_5194, n_5195, n_5196, n_5197, a_SCH2ADDRREG_F9_G_aCLRN, a_EQ1004,
          n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211,
          n_5212, a_SCH2ADDRREG_F9_G_aCLK, a_N2549, a_EQ606, n_5216, n_5217,
          n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225,
          n_5226, n_5227, n_5228, a_LC4_A8, a_EQ657, n_5231, n_5232, n_5233,
          n_5234, n_5235, n_5236, n_5237, n_5238, a_SCH0ADDRREG_F9_G, n_5240,
          n_5241, n_5242, n_5243, a_LC3_A8, a_EQ658, n_5246, n_5247, n_5248,
          n_5249, n_5250, n_5251, n_5252, n_5253, a_SCH0ADDRREG_F9_G_aCLRN,
          a_EQ876, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, n_5266,
          n_5267, n_5268, a_SCH0ADDRREG_F9_G_aCLK, a_LC2_A12, a_EQ683, n_5272,
          n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, a_SCH1ADDRREG_F9_G,
          n_5281, n_5282, n_5283, n_5284, a_LC3_A12, a_EQ684, n_5287, n_5288,
          n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, a_SCH1ADDRREG_F9_G_aCLRN,
          a_EQ940, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307,
          n_5308, n_5309, a_SCH1ADDRREG_F9_G_aCLK, a_LC2_A21, a_EQ824, n_5313,
          n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, a_SCH3WRDCNTREG_F9_G,
          n_5321, a_LC1_A21, a_EQ825, n_5324, n_5325, n_5326, n_5327, n_5328,
          n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, a_SCH3WRDCNTREG_F9_G_aCLRN,
          a_EQ1122, n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348,
          n_5349, n_5350, a_SCH3WRDCNTREG_F9_G_aCLK, a_N2367, a_EQ563, n_5354,
          n_5355, n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, n_5362,
          n_5363, a_N824, a_N824_aCLRN, a_N824_aD, n_5371, n_5372, n_5373,
          n_5375, n_5376, a_N824_aCLK, a_LC2_B15, a_LC2_B15_aIN, n_5380, n_5381,
          n_5382, n_5383, n_5384, n_5386, a_N2592, a_EQ643, n_5389, n_5390,
          n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398,
          a_N1523, a_EQ457, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406,
          a_STCSTATUS_F1_G, a_STCSTATUS_F1_G_aCLRN, a_EQ1178, n_5414, n_5415,
          n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423,
          a_STCSTATUS_F1_G_aCLK, a_LC5_C4, a_EQ831, n_5427, n_5428, n_5429,
          n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, a_N1047_aNOT,
          a_N1047_aNOT_aIN, n_5439, n_5440, n_5441, n_5442, n_5443, a_SCH3WRDCNTREG_F2_G_aCLRN,
          a_EQ1115, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456,
          n_5457, n_5458, n_5459, a_SCH3WRDCNTREG_F2_G_aCLK, a_LC1_D20, a_EQ811,
          n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470,
          n_5471, n_5472, a_N799, a_N799_aIN, n_5475, n_5476, n_5477, n_5478,
          n_5479, a_SCH2WRDCNTREG_F2_G_aCLRN, a_EQ1051, n_5486, n_5487, n_5488,
          n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, a_SCH2WRDCNTREG_F2_G_aCLK,
          a_LC3_C3, a_EQ769, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504,
          n_5505, n_5506, a_LC5_C3, a_EQ770, n_5509, n_5510, n_5511, n_5512,
          n_5513, n_5514, n_5515, n_5516, a_SCH0WRDCNTREG_F2_G_aCLRN, a_EQ923,
          n_5523, n_5524, n_5525, n_5526, n_5527, n_5528, n_5529, n_5530,
          n_5531, a_SCH0WRDCNTREG_F2_G_aCLK, a_LC3_D26, a_EQ792, n_5535, n_5536,
          n_5537, n_5538, n_5539, n_5540, a_SCH1BWORDOUT_F2_G, n_5542, n_5543,
          a_N434, a_N434_aIN, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551,
          n_5552, a_SCH1WRDCNTREG_F2_G_aCLRN, a_EQ987, n_5559, n_5560, n_5561,
          n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, a_SCH1WRDCNTREG_F2_G_aCLK,
          a_LC2_A9, a_EQ006, n_5572, n_5573, n_5574, n_5575, n_5576, a_SADDRESSOUT_F10_G,
          n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585,
          n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593,
          n_5594, n_5595, n_5596, n_5597, n_5598, a_LC3_E20, a_EQ709, n_5601,
          n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608, a_SCH2ADDRREG_F10_G,
          n_5610, n_5611, n_5612, n_5613, a_LC4_E20, a_EQ710, n_5616, n_5617,
          n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624, n_5625,
          n_5626, n_5627, n_5628, a_SCH2ADDRREG_F10_G_aCLRN, a_EQ1005, n_5635,
          n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642, n_5643,
          a_SCH2ADDRREG_F10_G_aCLK, a_LC4_E5, a_EQ822, n_5647, n_5648, n_5649,
          n_5650, n_5651, n_5652, n_5653, a_SH3WRDCNTREG_F10_G, n_5655, a_LC3_E5,
          a_EQ823, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664,
          n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, a_SH3WRDCNTREG_F10_G_aCLRN,
          a_EQ1151, n_5677, n_5678, n_5679, n_5680, n_5681, n_5682, n_5683,
          n_5684, n_5685, a_SH3WRDCNTREG_F10_G_aCLK, a_LC6_E9, a_EQ734, n_5689,
          n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696, a_SCH3ADDRREG_F10_G,
          n_5698, n_5699, n_5700, n_5701, a_LC4_E9, a_EQ735, n_5704, n_5705,
          n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713,
          n_5714, n_5715, n_5716, a_SCH3ADDRREG_F10_G_aCLRN, a_EQ1069, n_5723,
          n_5724, n_5725, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731,
          a_SCH3ADDRREG_F10_G_aCLK, a_LC1_E17, a_EQ801, n_5735, n_5736, n_5737,
          n_5738, n_5739, n_5740, n_5741, n_5742, a_SH2WRDCNTREG_F10_G, n_5744,
          n_5745, n_5746, n_5747, a_LC2_E17, a_EQ802, n_5750, n_5751, n_5752,
          n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760,
          n_5761, n_5762, a_SH2WRDCNTREG_F10_G_aCLRN, a_EQ1145, n_5769, n_5770,
          n_5771, n_5772, n_5773, n_5774, n_5775, n_5776, n_5777, a_SH2WRDCNTREG_F10_G_aCLK,
          a_N2550, a_EQ607, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786,
          n_5787, n_5788, n_5789, n_5790, n_5791, n_5792, n_5793, a_LC4_E11,
          a_EQ681, n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802,
          n_5803, a_SCH1ADDRREG_F10_G, n_5805, n_5806, n_5807, n_5808, a_LC5_E11,
          a_EQ682, n_5811, n_5812, n_5813, n_5814, n_5815, n_5816, n_5817,
          n_5818, a_SCH1ADDRREG_F10_G_aCLRN, a_EQ941, n_5825, n_5826, n_5827,
          n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, a_SCH1ADDRREG_F10_G_aCLK,
          a_LC6_E17, a_EQ222, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842,
          n_5843, n_5844, a_SH0WRDCNTREG_F10_G, n_5846, n_5847, n_5848, n_5849,
          a_LC3_E17, a_EQ221, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857,
          n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, a_SH0WRDCNTREG_F10_G_aCLRN,
          a_EQ1133, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877,
          n_5878, n_5879, a_SH0WRDCNTREG_F10_G_aCLK, a_LC4_E13, a_EQ655, n_5883,
          n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, a_SCH0ADDRREG_F10_G,
          n_5892, n_5893, n_5894, n_5895, a_LC5_E13, a_EQ656, n_5898, n_5899,
          n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, a_SCH0ADDRREG_F10_G_aCLRN,
          a_EQ877, n_5912, n_5913, n_5914, n_5915, n_5916, n_5917, n_5918,
          n_5919, n_5920, a_SCH0ADDRREG_F10_G_aCLK, a_LC3_E12, a_EQ780, n_5924,
          n_5925, n_5926, n_5927, a_SH1WRDCNTREG_F10_G, n_5929, n_5930, a_SCH1BWORDOUT_F10_G,
          n_5932, n_5933, a_LC4_E12, a_EQ781, n_5936, n_5937, n_5938, n_5939,
          n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947,
          a_SH1WRDCNTREG_F10_G_aCLRN, a_EQ1139, n_5954, n_5955, n_5956, n_5957,
          n_5958, n_5959, n_5960, n_5961, n_5962, a_SH1WRDCNTREG_F10_G_aCLK,
          a_LC3_A9, a_EQ013, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971,
          n_5972, n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979,
          n_5980, a_LC8_A9, a_EQ007, n_5983, n_5984, n_5985, n_5986, a_SADDRESSOUT_F11_G,
          n_5988, n_5989, n_5990, n_5991, a_LC1_A16, a_EQ707, n_5994, n_5995,
          n_5996, n_5997, n_5998, n_5999, n_6000, a_SCH2ADDRREG_F11_G, n_6002,
          a_LC2_A16, a_EQ708, n_6005, n_6006, n_6007, n_6008, n_6009, n_6010,
          n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, a_SCH2ADDRREG_F11_G_aCLRN,
          a_EQ1006, n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030,
          n_6031, n_6032, a_SCH2ADDRREG_F11_G_aCLK, a_LC5_F1, a_EQ732, n_6036,
          n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, a_SCH3ADDRREG_F11_G,
          n_6045, n_6046, n_6047, n_6048, a_LC2_F1, a_EQ733, n_6051, n_6052,
          n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060,
          n_6061, n_6062, n_6063, a_SCH3ADDRREG_F11_G_aCLRN, a_EQ1070, n_6070,
          n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078,
          a_SCH3ADDRREG_F11_G_aCLK, a_N2551, a_EQ608, n_6082, n_6083, n_6084,
          n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092,
          n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100,
          n_6101, n_6102, n_6103, n_6104, a_LC4_A24, a_EQ653, n_6107, n_6108,
          n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, a_SCH0ADDRREG_F11_G,
          n_6116, n_6117, n_6118, n_6119, a_LC6_A24, a_EQ654, n_6122, n_6123,
          n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, a_SCH0ADDRREG_F11_G_aCLRN,
          a_EQ878, n_6136, n_6137, n_6138, n_6139, n_6140, n_6141, n_6142,
          n_6143, n_6144, a_SCH0ADDRREG_F11_G_aCLK, a_LC1_A23, a_EQ679, n_6148,
          n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6155, a_SCH1ADDRREG_F11_G,
          n_6157, n_6158, n_6159, n_6160, a_LC2_A23, a_EQ680, n_6163, n_6164,
          n_6165, n_6166, n_6167, n_6168, n_6169, n_6170, a_SCH1ADDRREG_F11_G_aCLRN,
          a_EQ942, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183,
          n_6184, n_6185, a_SCH1ADDRREG_F11_G_aCLK, a_LC4_C20, a_EQ830, n_6189,
          n_6190, n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197,
          n_6198, a_N1036_aNOT, a_N1036_aNOT_aIN, n_6201, n_6202, n_6203,
          n_6204, n_6205, a_SCH3WRDCNTREG_F3_G_aCLRN, a_EQ1116, n_6212, n_6213,
          n_6214, n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221,
          a_SCH3WRDCNTREG_F3_G_aCLK, a_LC5_A9, a_EQ008, n_6225, n_6226, n_6227,
          n_6228, n_6229, a_SADDRESSOUT_F12_G, n_6231, n_6232, n_6233, n_6234,
          n_6235, n_6236, n_6237, n_6238, n_6239, n_6240, n_6241, n_6242,
          n_6243, n_6244, n_6245, n_6246, n_6247, n_6248, n_6249, n_6250,
          n_6251, a_LC4_A14, a_EQ705, n_6254, n_6255, n_6256, n_6257, n_6258,
          n_6259, n_6260, a_SCH2ADDRREG_F12_G, n_6262, a_LC5_A14, a_EQ706,
          n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271, n_6272,
          n_6273, n_6274, n_6275, n_6276, n_6277, a_SCH2ADDRREG_F12_G_aCLRN,
          a_EQ1007, n_6284, n_6285, n_6286, n_6287, n_6288, n_6289, n_6290,
          n_6291, n_6292, a_SCH2ADDRREG_F12_G_aCLK, a_N2552, a_EQ609, n_6296,
          n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303, n_6304,
          n_6305, n_6306, n_6307, n_6308, a_N212, a_N212_aIN, n_6311, n_6312,
          n_6313, n_6314, n_6315, a_N217, a_EQ213, n_6318, n_6319, n_6320,
          n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, a_SCH0ADDRREG_F12_G,
          n_6328, a_SCH0ADDRREG_F12_G_aCLRN, a_EQ879, n_6335, n_6336, n_6337,
          n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344, n_6345,
          n_6346, a_SCH0ADDRREG_F12_G_aCLK, a_LC2_A15, a_EQ730, n_6350, n_6351,
          n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, a_SCH3ADDRREG_F12_G,
          n_6359, n_6360, n_6361, n_6362, a_LC1_A15, a_EQ731, n_6365, n_6366,
          n_6367, n_6368, n_6369, n_6370, n_6371, n_6372, n_6373, n_6374,
          n_6375, n_6376, n_6377, a_SCH3ADDRREG_F12_G_aCLRN, a_EQ1071, n_6384,
          n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392,
          a_SCH3ADDRREG_F12_G_aCLK, a_LC3_F18, a_LC3_F18_aIN, n_6396, n_6397,
          n_6398, n_6399, n_6400, n_6401, a_LC8_A12, a_EQ678, n_6404, n_6405,
          n_6406, n_6407, a_SCH1ADDRREG_F12_G, n_6409, n_6410, n_6411, n_6412,
          a_N443, a_N443_aIN, n_6415, n_6416, n_6417, n_6418, n_6419, n_6420,
          n_6421, a_SCH1ADDRREG_F12_G_aCLRN, a_EQ943, n_6428, n_6429, n_6430,
          n_6431, n_6432, n_6433, n_6434, n_6435, n_6436, n_6437, a_SCH1ADDRREG_F12_G_aCLK,
          a_N66, a_N66_aIN, n_6441, n_6442, n_6443, n_6444, n_6445, n_6446,
          n_6447, a_N2569_aNOT, a_EQ622, n_6450, n_6451, n_6452, n_6453, n_6454,
          n_6455, n_6456, n_6457, n_6458, n_6459, a_SCH2MODEREG_F3_G_aCLRN,
          a_EQ1046, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472,
          n_6473, n_6474, a_SCH2MODEREG_F3_G_aCLK, a_N2532_aNOT, a_N2532_aNOT_aIN,
          n_6478, n_6479, n_6480, n_6481, n_6482, a_N2567, a_N2567_aIN, n_6485,
          n_6486, n_6487, n_6488, n_6489, n_6490, a_SCH0MODEREG_F3_G_aCLRN,
          a_EQ918, n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503,
          n_6504, n_6505, a_SCH0MODEREG_F3_G_aCLK, a_N84, a_N84_aIN, n_6509,
          n_6510, n_6511, n_6512, n_6513, a_N2568, a_N2568_aIN, n_6516, n_6517,
          n_6518, n_6519, n_6520, n_6521, a_SCH1MODEREG_F3_G_aCLRN, a_EQ982,
          n_6528, n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535,
          n_6536, a_SCH1MODEREG_F3_G_aCLK, a_N2570_aNOT, a_EQ623, n_6540,
          n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548,
          n_6549, a_SCH3MODEREG_F3_G_aCLRN, a_EQ1110, n_6556, n_6557, n_6558,
          n_6559, n_6560, n_6561, n_6562, n_6563, n_6564, a_SCH3MODEREG_F3_G_aCLK,
          a_LC5_F8, a_EQ263, n_6568, n_6569, n_6570, n_6571, n_6572, n_6573,
          n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580, n_6581,
          n_6582, a_LC6_F8, a_EQ764, n_6585, n_6586, n_6587, n_6588, n_6589,
          n_6590, n_6591, n_6592, n_6593, n_6594, a_SCH0WRDCNTREG_F5_G_aCLRN,
          a_EQ926, n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607,
          n_6608, n_6609, n_6610, n_6611, n_6612, a_SCH0WRDCNTREG_F5_G_aCLK,
          a_LC8_F2, a_EQ828, n_6616, n_6617, n_6618, n_6619, n_6620, n_6621,
          n_6622, n_6623, n_6624, n_6625, a_N1061_aNOT, a_EQ348, n_6628, n_6629,
          n_6630, n_6631, n_6632, n_6633, n_6634, n_6635, n_6636, n_6637,
          n_6638, n_6639, n_6640, n_6641, n_6642, a_SCH3WRDCNTREG_F5_G_aCLRN,
          a_EQ1118, n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655,
          n_6656, n_6657, n_6658, a_SCH3WRDCNTREG_F5_G_aCLK, a_LC3_F2, a_EQ252,
          n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668, n_6669,
          n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676, a_LC4_F2,
          a_EQ787, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684, n_6685,
          n_6686, n_6687, n_6688, a_SCH1WRDCNTREG_F5_G_aCLRN, a_EQ990, n_6695,
          n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703,
          n_6704, n_6705, n_6706, a_SCH1WRDCNTREG_F5_G_aCLK, a_LC6_F24, a_EQ808,
          n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716, n_6717,
          n_6718, n_6719, a_N833_aNOT, a_EQ312, n_6722, n_6723, n_6724, n_6725,
          n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732, n_6733,
          n_6734, n_6735, n_6736, a_SCH2WRDCNTREG_F5_G_aCLRN, a_EQ1054, n_6743,
          n_6744, n_6745, n_6746, n_6747, n_6748, n_6749, n_6750, n_6751,
          n_6752, a_SCH2WRDCNTREG_F5_G_aCLK, a_LC1_E6, a_EQ752, n_6756, n_6757,
          n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, a_SH0WRDCNTREG_F13_G,
          n_6765, n_6766, n_6767, n_6768, a_LC2_E6, a_EQ753, n_6771, n_6772,
          n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780,
          n_6781, n_6782, n_6783, a_SH0WRDCNTREG_F13_G_aCLRN, a_EQ1136, n_6790,
          n_6791, n_6792, n_6793, n_6794, n_6795, n_6796, n_6797, n_6798,
          a_SH0WRDCNTREG_F13_G_aCLK, a_LC3_E25, a_EQ816, n_6802, n_6803, n_6804,
          n_6805, n_6806, n_6807, n_6808, a_SH3WRDCNTREG_F13_G, n_6810, a_LC4_E25,
          a_EQ817, n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819,
          n_6820, n_6821, n_6822, n_6823, n_6824, n_6825, a_SH3WRDCNTREG_F13_G_aCLRN,
          a_EQ1154, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837, n_6838,
          n_6839, n_6840, a_SH3WRDCNTREG_F13_G_aCLK, a_LC1_E19, a_EQ774, n_6844,
          n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, a_SH1WRDCNTREG_F13_G,
          n_6852, a_LC4_E19, a_EQ775, n_6855, n_6856, n_6857, n_6858, n_6859,
          n_6860, n_6861, n_6862, n_6863, n_6864, n_6865, n_6866, n_6867,
          a_SH1WRDCNTREG_F13_G_aCLRN, a_EQ1142, n_6874, n_6875, n_6876, n_6877,
          n_6878, n_6879, n_6880, n_6881, n_6882, a_SH1WRDCNTREG_F13_G_aCLK,
          a_LC1_A9, a_EQ012, n_6886, n_6887, n_6888, n_6889, n_6890, n_6891,
          n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6898, n_6899,
          n_6900, a_N2594_aNOT, a_EQ644, n_6903, n_6904, n_6905, n_6906, n_6907,
          a_SADDRESSOUT_F13_G, n_6909, n_6910, n_6911, n_6912, n_6913, n_6914,
          n_6915, n_6916, n_6917, n_6918, n_6919, n_6920, n_6921, n_6922,
          n_6923, n_6924, n_6925, n_6926, a_LC7_F25, a_EQ677, n_6929, n_6930,
          n_6931, n_6932, a_SCH1ADDRREG_F13_G, n_6934, n_6935, n_6936, n_6937,
          a_N436, a_N436_aIN, n_6940, n_6941, n_6942, n_6943, n_6944, n_6945,
          n_6946, a_SCH1ADDRREG_F13_G_aCLRN, a_EQ944, n_6953, n_6954, n_6955,
          n_6956, n_6957, n_6958, n_6959, n_6960, n_6961, n_6962, a_SCH1ADDRREG_F13_G_aCLK,
          a_LC5_E25, a_EQ795, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971,
          n_6972, n_6973, a_SH2WRDCNTREG_F13_G, n_6975, n_6976, n_6977, n_6978,
          a_LC6_E25, a_EQ796, n_6981, n_6982, n_6983, n_6984, n_6985, n_6986,
          n_6987, n_6988, n_6989, n_6990, n_6991, n_6992, n_6993, a_SH2WRDCNTREG_F13_G_aCLRN,
          a_EQ1148, n_7000, n_7001, n_7002, n_7003, n_7004, n_7005, n_7006,
          n_7007, n_7008, a_SH2WRDCNTREG_F13_G_aCLK, a_LC7_E3, a_EQ009, n_7012,
          n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, a_LC1_E20,
          a_EQ703, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028,
          a_SCH2ADDRREG_F13_G, n_7030, a_LC2_E20, a_EQ704, n_7033, n_7034,
          n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041, n_7042,
          n_7043, n_7044, n_7045, a_SCH2ADDRREG_F13_G_aCLRN, a_EQ1008, n_7052,
          n_7053, n_7054, n_7055, n_7056, n_7057, n_7058, n_7059, n_7060,
          a_SCH2ADDRREG_F13_G_aCLK, a_N218, a_EQ214, n_7064, n_7065, n_7066,
          n_7067, n_7068, n_7069, n_7070, a_SCH0ADDRREG_F13_G, n_7072, n_7073,
          n_7074, a_N216, a_EQ212, n_7077, n_7078, n_7079, n_7080, n_7081,
          n_7082, a_SCH0ADDRREG_F13_G_aCLRN, a_EQ880, n_7089, n_7090, n_7091,
          n_7092, n_7093, n_7094, n_7095, n_7096, n_7097, n_7098, a_SCH0ADDRREG_F13_G_aCLK,
          a_LC2_E9, a_EQ728, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107,
          n_7108, n_7109, a_SCH3ADDRREG_F13_G, n_7111, n_7112, n_7113, n_7114,
          a_LC1_E9, a_EQ729, n_7117, n_7118, n_7119, n_7120, n_7121, n_7122,
          n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129, a_SCH3ADDRREG_F13_G_aCLRN,
          a_EQ1072, n_7136, n_7137, n_7138, n_7139, n_7140, n_7141, n_7142,
          n_7143, n_7144, a_SCH3ADDRREG_F13_G_aCLK, a_SCH1MODEREG_F4_G, a_SCH1MODEREG_F4_G_aCLRN,
          a_EQ983, n_7153, n_7154, n_7155, n_7156, n_7157, n_7158, n_7159,
          n_7160, n_7161, a_SCH1MODEREG_F4_G_aCLK, a_SCH2MODEREG_F4_G, a_SCH2MODEREG_F4_G_aCLRN,
          a_EQ1047, n_7170, n_7171, n_7172, n_7173, n_7174, n_7175, n_7176,
          n_7177, n_7178, a_SCH2MODEREG_F4_G_aCLK, a_SCH3MODEREG_F4_G, a_SCH3MODEREG_F4_G_aCLRN,
          a_EQ1111, n_7187, n_7188, n_7189, n_7190, n_7191, n_7192, n_7193,
          n_7194, n_7195, a_SCH3MODEREG_F4_G_aCLK, a_SCH0MODEREG_F4_G, a_SCH0MODEREG_F4_G_aCLRN,
          a_EQ919, n_7204, n_7205, n_7206, n_7207, n_7208, n_7209, n_7210,
          n_7211, n_7212, a_SCH0MODEREG_F4_G_aCLK, a_LC6_F12, a_EQ011, n_7216,
          n_7217, n_7218, n_7219, n_7220, n_7221, n_7222, n_7223, n_7224,
          n_7225, n_7226, n_7227, n_7228, a_LC1_F12, a_EQ010, n_7231, n_7232,
          n_7233, n_7234, a_SADDRESSOUT_F14_G, n_7236, n_7237, n_7238, n_7239,
          a_N2554, a_EQ610, n_7242, n_7243, n_7244, n_7245, n_7246, n_7247,
          n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7254, a_LC3_F7,
          a_EQ651, n_7257, n_7258, n_7259, n_7260, n_7261, n_7262, n_7263,
          a_SCH0ADDRREG_F14_G, n_7265, a_LC4_F7, a_EQ652, n_7268, n_7269,
          n_7270, n_7271, n_7272, n_7273, n_7274, n_7275, a_SCH0ADDRREG_F14_G_aCLRN,
          a_EQ881, n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288,
          n_7289, n_7290, a_SCH0ADDRREG_F14_G_aCLK, a_LC1_F22, a_EQ701, n_7294,
          n_7295, n_7296, n_7297, n_7298, n_7299, n_7300, a_SCH2ADDRREG_F14_G,
          n_7302, a_LC3_F22, a_EQ702, n_7305, n_7306, n_7307, n_7308, n_7309,
          n_7310, n_7311, n_7312, a_SCH2ADDRREG_F14_G_aCLRN, a_EQ1009, n_7319,
          n_7320, n_7321, n_7322, n_7323, n_7324, n_7325, n_7326, n_7327,
          n_7328, n_7329, n_7330, n_7331, a_SCH2ADDRREG_F14_G_aCLK, a_LC8_F25,
          a_EQ676, n_7335, n_7336, n_7337, n_7338, a_SCH1ADDRREG_F14_G, n_7340,
          n_7341, n_7342, n_7343, a_N440, a_N440_aIN, n_7346, n_7347, n_7348,
          n_7349, n_7350, n_7351, n_7352, a_SCH1ADDRREG_F14_G_aCLRN, a_EQ945,
          n_7359, n_7360, n_7361, n_7362, n_7363, n_7364, n_7365, n_7366,
          n_7367, n_7368, a_SCH1ADDRREG_F14_G_aCLK, a_LC4_F1, a_EQ726, n_7372,
          n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, a_SCH3ADDRREG_F14_G,
          n_7381, n_7382, n_7383, n_7384, a_LC3_F1, a_EQ727, n_7387, n_7388,
          n_7389, n_7390, n_7391, n_7392, n_7393, n_7394, n_7395, n_7396,
          n_7397, n_7398, n_7399, a_SCH3ADDRREG_F14_G_aCLRN, a_EQ1073, n_7406,
          n_7407, n_7408, n_7409, n_7410, n_7411, n_7412, n_7413, n_7414,
          a_SCH3ADDRREG_F14_G_aCLK, a_LC4_D2, a_EQ826, n_7418, n_7419, n_7420,
          n_7421, n_7422, n_7423, n_7424, n_7425, n_7426, a_SCH3WRDCNTREG_F7_G,
          n_7428, a_N1038_aNOT, a_EQ345, n_7431, n_7432, n_7433, n_7434, n_7435,
          n_7436, n_7437, n_7438, n_7439, n_7440, a_SCH3WRDCNTREG_F7_G_aCLRN,
          a_EQ1120, n_7447, n_7448, n_7449, n_7450, n_7451, n_7452, n_7453,
          n_7454, n_7455, n_7456, a_SCH3WRDCNTREG_F7_G_aCLK, a_N782_aNOT,
          a_EQ298, n_7460, n_7461, n_7462, n_7463, n_7464, n_7465, n_7466,
          a_SCH2WRDCNTREG_F7_G, n_7468, a_LC5_D5, a_EQ806, n_7471, n_7472,
          n_7473, n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480,
          n_7481, n_7482, n_7483, a_SCH2WRDCNTREG_F7_G_aCLRN, a_EQ1056, n_7490,
          n_7491, n_7492, n_7493, n_7494, n_7495, n_7496, n_7497, n_7498,
          a_SCH2WRDCNTREG_F7_G_aCLK, a_N646_aNOT, a_EQ278, n_7502, n_7503,
          n_7504, n_7505, n_7506, n_7507, n_7508, a_SCH1WRDCNTREG_F7_G, n_7510,
          a_LC4_D11, a_EQ784, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518,
          n_7519, n_7520, n_7521, a_SCH1WRDCNTREG_F7_G_aCLRN, a_EQ992, n_7528,
          n_7529, n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536,
          n_7537, n_7538, n_7539, n_7540, a_SCH1WRDCNTREG_F7_G_aCLK, a_LC4_D9,
          a_EQ760, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550,
          a_SCH0WRDCNTREG_F7_G, n_7552, a_LC5_D9, a_EQ761, n_7555, n_7556,
          n_7557, n_7558, n_7559, n_7560, n_7561, n_7562, n_7563, n_7564,
          n_7565, n_7566, n_7567, a_SCH0WRDCNTREG_F7_G_aCLRN, a_EQ928, n_7574,
          n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581, n_7582,
          a_SCH0WRDCNTREG_F7_G_aCLK, a_LC3_F12, a_EQ834, n_7586, n_7587, n_7588,
          n_7589, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596,
          n_7597, n_7598, n_7599, a_N3045, a_EQ835, n_7602, n_7603, n_7604,
          n_7605, a_SADDRESSOUT_F15_G, n_7607, n_7608, n_7609, n_7610, a_LC6_D5,
          a_EQ700, n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619,
          n_7620, a_SCH2ADDRREG_F15_G, n_7622, a_N818, a_N818_aIN, n_7625,
          n_7626, n_7627, n_7628, n_7629, n_7630, a_SCH2ADDRREG_F15_G_aCLRN,
          a_EQ1010, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643,
          n_7644, n_7645, n_7646, n_7647, a_SCH2ADDRREG_F15_G_aCLK, a_N2555,
          a_EQ611, n_7651, n_7652, n_7653, n_7654, n_7655, n_7656, n_7657,
          n_7658, a_LC2_D10, a_EQ649, n_7661, n_7662, n_7663, n_7664, n_7665,
          n_7666, n_7667, n_7668, a_SCH0ADDRREG_F15_G, n_7670, n_7671, n_7672,
          n_7673, a_LC1_D10, a_EQ650, n_7676, n_7677, n_7678, n_7679, n_7680,
          n_7681, n_7682, n_7683, a_SCH0ADDRREG_F15_G_aCLRN, a_EQ882, n_7690,
          n_7691, n_7692, n_7693, n_7694, n_7695, n_7696, n_7697, n_7698,
          a_SCH0ADDRREG_F15_G_aCLK, a_LC6_D3, a_EQ724, n_7702, n_7703, n_7704,
          n_7705, n_7706, n_7707, n_7708, n_7709, a_SCH3ADDRREG_F15_G, n_7711,
          n_7712, n_7713, n_7714, a_LC5_D3, a_EQ725, n_7717, n_7718, n_7719,
          n_7720, n_7721, n_7722, n_7723, n_7724, a_SCH3ADDRREG_F15_G_aCLRN,
          a_EQ1074, n_7731, n_7732, n_7733, n_7734, n_7735, n_7736, n_7737,
          n_7738, n_7739, a_SCH3ADDRREG_F15_G_aCLK, a_LC5_D11, a_EQ675, n_7743,
          n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750, a_SCH1ADDRREG_F15_G,
          n_7752, a_N457, a_N457_aIN, n_7755, n_7756, n_7757, n_7758, n_7759,
          n_7760, n_7761, a_SCH1ADDRREG_F15_G_aCLRN, a_EQ946, n_7768, n_7769,
          n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776, n_7777,
          n_7778, a_SCH1ADDRREG_F15_G_aCLK, a_N63_aNOT, a_EQ184, n_7782, n_7783,
          n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790, n_7791,
          a_N2566_aNOT, a_EQ619, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799,
          a_N1434_aNOT, a_EQ439, n_7802, n_7803, n_7804, n_7805, n_7806, a_SREQUESTREG_F1_G,
          n_7808, n_7809, n_7810, n_7811, n_7812, a_SREQUESTREG_F1_G_aCLRN,
          a_EQ1174, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824, n_7825,
          n_7826, n_7827, a_SREQUESTREG_F1_G_aCLK, a_N2582_aNOT, a_EQ634,
          n_7831, n_7832, n_7833, n_7834, n_7835, n_7836, a_SCH2BAROUT_F1_G,
          a_SCH2BAROUT_F1_G_aCLRN, a_EQ1012, n_7844, n_7845, n_7846, n_7847,
          n_7848, n_7849, n_7850, n_7851, n_7852, a_SCH2BAROUT_F1_G_aCLK,
          a_N2580_aNOT, a_EQ631, n_7856, n_7857, n_7858, n_7859, n_7860, n_7861,
          a_SCH3BAROUT_F5_G, a_SCH3BAROUT_F5_G_aCLRN, a_EQ1080, n_7869, n_7870,
          n_7871, n_7872, n_7873, n_7874, n_7875, n_7876, n_7877, a_SCH3BAROUT_F5_G_aCLK,
          a_SCH3BAROUT_F7_G, a_SCH3BAROUT_F7_G_aCLRN, a_EQ1082, n_7886, n_7887,
          n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, a_SCH3BAROUT_F7_G_aCLK,
          a_LC3_D21, a_EQ748, n_7898, n_7899, n_7900, n_7901, n_7902, n_7903,
          n_7904, n_7905, a_SH0WRDCNTREG_F15_G, n_7907, n_7908, n_7909, n_7910,
          a_LC5_D21, a_EQ749, n_7913, n_7914, n_7915, n_7916, n_7917, n_7918,
          n_7919, n_7920, n_7921, n_7922, n_7923, n_7924, n_7925, a_SH0WRDCNTREG_F15_G_aCLRN,
          a_EQ1138, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937, n_7938,
          n_7939, n_7940, a_SH0WRDCNTREG_F15_G_aCLK, a_LC7_D4, a_EQ315, n_7944,
          n_7945, n_7946, n_7947, n_7948, n_7949, n_7950, a_SH1WRDCNTREG_F15_G,
          n_7952, a_LC5_D4, a_EQ324, n_7955, n_7956, n_7957, n_7958, n_7959,
          n_7960, n_7961, n_7962, n_7963, n_7964, n_7965, n_7966, n_7967,
          a_SH1WRDCNTREG_F15_G_aCLRN, a_EQ1144, n_7974, n_7975, n_7976, n_7977,
          n_7978, n_7979, n_7980, n_7981, n_7982, a_SH1WRDCNTREG_F15_G_aCLK,
          a_N1149_aNOT, a_EQ370, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991,
          n_7992, n_7993, a_SH2WRDCNTREG_F15_G, n_7995, n_7996, n_7997, n_7998,
          a_LC1_D7, a_EQ371, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006,
          n_8007, n_8008, n_8009, n_8010, n_8011, n_8012, n_8013, a_SH2WRDCNTREG_F15_G_aCLRN,
          a_EQ1150, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025, n_8026,
          n_8027, n_8028, a_SH2WRDCNTREG_F15_G_aCLK, a_LC2_D3, a_EQ814, n_8032,
          n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, a_SH3WRDCNTREG_F15_G,
          n_8040, a_LC3_D3, a_EQ815, n_8043, n_8044, n_8045, n_8046, n_8047,
          n_8048, n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055,
          a_SH3WRDCNTREG_F15_G_aCLRN, a_EQ1156, n_8062, n_8063, n_8064, n_8065,
          n_8066, n_8067, n_8068, n_8069, n_8070, a_SH3WRDCNTREG_F15_G_aCLK,
          a_LC2_D24, a_EQ277, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079,
          n_8080, n_8081, n_8082, n_8083, n_8084, n_8085, a_LC4_D24, a_EQ276,
          n_8088, n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095,
          a_N629_aNOT, a_EQ274, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103,
          n_8104, n_8105, a_LC4_D15, a_EQ273, n_8108, n_8109, n_8110, n_8111,
          n_8112, n_8113, n_8114, n_8115, a_LC2_D15, a_EQ272, n_8118, n_8119,
          n_8120, n_8121, n_8122, n_8123, n_8124, n_8125, a_N3549_aCLRN, a_EQ845,
          n_8132, n_8133, n_8134, n_8135, n_8136, n_8137, n_8138, n_8139,
          n_8140, n_8141, n_8142, n_8143, a_N3549_aCLK, a_N1174, a_EQ381,
          n_8147, n_8148, n_8149, n_8150, n_8151, n_8152, n_8153, n_8154,
          a_N1163_aNOT, a_EQ373, n_8157, n_8158, n_8159, n_8160, n_8161, n_8162,
          n_8163, n_8164, a_LC6_D24, a_EQ382, n_8167, n_8168, n_8169, n_8170,
          n_8171, n_8172, n_8173, n_8174, a_LC1_D6, a_EQ380, n_8177, n_8178,
          n_8179, n_8180, n_8181, n_8182, n_8183, n_8184, a_LC1_D24, a_EQ379,
          n_8187, n_8188, n_8189, n_8190, n_8191, n_8192, n_8193, n_8194,
          a_N3548_aCLRN, a_EQ844, n_8201, n_8202, n_8203, n_8204, n_8205,
          n_8206, n_8207, n_8208, n_8209, n_8210, n_8211, n_8212, a_N3548_aCLK,
          a_LC5_A13, a_EQ227, n_8216, n_8217, n_8218, n_8219, n_8220, n_8221,
          n_8222, n_8223, a_LC2_A13, a_EQ225, n_8226, n_8227, n_8228, n_8229,
          n_8230, n_8231, n_8232, n_8233, n_8234, n_8235, n_8236, a_N295_aNOT,
          a_EQ226, n_8239, n_8240, n_8241, n_8242, n_8243, n_8244, n_8245,
          n_8246, a_LC8_A13, a_EQ229, n_8249, n_8250, n_8251, n_8252, n_8253,
          n_8254, n_8255, n_8256, a_LC7_A13, a_EQ228, n_8259, n_8260, n_8261,
          n_8262, n_8263, n_8264, n_8265, n_8266, a_N3547_aCLRN, a_EQ843,
          n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280,
          n_8281, n_8282, n_8283, n_8284, a_N3547_aCLK, a_N73, a_N73_aIN,
          n_8288, n_8289, n_8290, n_8291, n_8292, n_8293, n_8294, a_N65, a_N65_aIN,
          n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, a_N1119_aNOT,
          a_EQ359, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312,
          a_N1103_aNOT, a_EQ354, n_8315, n_8316, n_8317, n_8318, n_8319, a_SMASKREG_F0_G_aNOT,
          n_8321, n_8322, n_8323, n_8324, n_8325, a_N2564, a_N2564_aIN, n_8328,
          n_8329, n_8330, n_8331, n_8332, a_LC2_B4_aNOT, a_EQ356, n_8335,
          n_8336, n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343,
          a_N75_aNOT, a_EQ193, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351,
          n_8352, n_8353, n_8354, n_8355, a_N103_aNOT, a_N103_aNOT_aIN, n_8358,
          n_8359, n_8360, n_8361, n_8362, a_LC1_B4, a_EQ357, n_8365, n_8366,
          n_8367, n_8368, n_8369, n_8370, n_8371, a_N104_aNOT, a_N104_aNOT_aIN,
          n_8374, n_8375, n_8376, n_8377, n_8378, a_LC7_B4, a_EQ358, n_8381,
          n_8382, n_8383, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389,
          a_LC5_B4_aNOT, a_EQ353, n_8392, n_8393, n_8394, n_8395, n_8396,
          n_8397, n_8398, n_8399, a_N1108, a_EQ355, n_8402, n_8403, n_8404,
          n_8405, n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412,
          n_8413, a_N2565, a_N2565_aIN, n_8416, n_8417, n_8418, n_8419, n_8420,
          a_SMASKREG_F0_G_aNOT_aCLRN, a_EQ1157, n_8427, n_8428, n_8429, n_8430,
          n_8431, n_8432, n_8433, n_8434, n_8435, n_8436, a_SMASKREG_F0_G_aNOT_aCLK,
          a_N45, a_N45_aIN, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445,
          a_SREQUESTREG_F0_G, a_SREQUESTREG_F0_G_aCLRN, a_EQ1173, n_8453,
          n_8454, n_8455, n_8456, n_8457, n_8458, n_8459, n_8460, n_8461,
          n_8462, n_8463, a_SREQUESTREG_F0_G_aCLK, a_N1530_aNOT, a_EQ458,
          n_8467, n_8468, n_8469, a_STCSTATUS_F0_G, n_8471, n_8472, n_8473,
          n_8474, n_8475, a_STCSTATUS_F0_G_aCLRN, a_EQ1177, n_8482, n_8483,
          n_8484, n_8485, n_8486, n_8487, n_8488, n_8489, n_8490, n_8491,
          n_8492, a_STCSTATUS_F0_G_aCLK, a_N1446, a_EQ445, n_8496, n_8497,
          n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, a_LC2_B22_aNOT,
          a_EQ441, n_8506, n_8507, n_8508, n_8509, n_8510, a_SMASKREG_F1_G_aNOT,
          n_8512, n_8513, n_8514, n_8515, n_8516, a_LC4_B19, a_EQ539, n_8519,
          n_8520, n_8521, n_8522, n_8523, n_8524, n_8525, n_8526, n_8527,
          a_LC1_B17, a_LC1_B17_aIN, n_8530, n_8531, n_8532, n_8533, n_8534,
          n_8535, n_8536, a_LC2_B17_aNOT, a_EQ444, n_8539, n_8540, n_8541,
          n_8542, n_8543, n_8544, n_8545, n_8546, n_8547, n_8548, n_8549,
          a_LC7_B17_aNOT, a_EQ446, n_8552, n_8553, n_8554, n_8555, n_8556,
          n_8557, n_8558, n_8559, n_8560, n_8561, a_LC6_B17_aNOT, a_EQ440,
          n_8564, n_8565, n_8566, n_8567, n_8568, n_8569, n_8570, n_8571,
          a_LC8_B17_aNOT, a_EQ540, n_8574, n_8575, n_8576, n_8577, n_8578,
          n_8579, n_8580, n_8581, n_8582, a_N1432, a_N1432_aIN, n_8585, n_8586,
          n_8587, n_8588, n_8589, a_N1442_aNOT, a_EQ442, n_8592, n_8593, n_8594,
          n_8595, n_8596, n_8597, n_8598, n_8599, n_8600, n_8601, a_SMASKREG_F1_G_aNOT_aCLRN,
          a_EQ1158, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613, n_8614,
          n_8615, a_SMASKREG_F1_G_aNOT_aCLK, a_LC4_B9_aNOT, a_LC4_B9_aNOT_aIN,
          n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8625, a_SREQUESTREG_F2_G,
          a_SREQUESTREG_F2_G_aCLRN, a_EQ1175, n_8633, n_8634, n_8635, n_8636,
          n_8637, n_8638, n_8639, n_8640, n_8641, n_8642, n_8643, a_SREQUESTREG_F2_G_aCLK,
          a_STCSTATUS_F2_G, a_STCSTATUS_F2_G_aCLRN, a_EQ1179, n_8652, n_8653,
          n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8660, n_8661,
          a_STCSTATUS_F2_G_aCLK, a_LC3_B19_aNOT, a_LC3_B19_aNOT_aIN, n_8665,
          n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, a_LC7_B19, a_EQ536,
          n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681,
          n_8682, n_8683, a_LC2_B19, a_EQ435, n_8686, n_8687, n_8688, n_8689,
          n_8690, a_SMASKREG_F2_G_aNOT, n_8692, n_8693, n_8694, n_8695, n_8696,
          a_LC6_B19, a_EQ537, n_8699, n_8700, n_8701, n_8702, n_8703, n_8704,
          n_8705, n_8706, n_8707, n_8708, a_N46, a_N46_aIN, n_8711, n_8712,
          n_8713, n_8714, n_8715, a_LC6_B22_aNOT, a_EQ535, n_8718, n_8719,
          n_8720, n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727,
          n_8728, a_LC5_B22_aNOT, a_EQ538, n_8731, n_8732, n_8733, n_8734,
          n_8735, n_8736, n_8737, n_8738, n_8739, a_LC8_B22_aNOT, a_EQ436,
          n_8742, n_8743, n_8744, n_8745, n_8746, n_8747, n_8748, n_8749,
          n_8750, n_8751, a_LC7_B22_aNOT, a_EQ534, n_8754, n_8755, n_8756,
          n_8757, n_8758, n_8759, n_8760, n_8761, a_SMASKREG_F2_G_aNOT_aCLRN,
          a_EQ1159, n_8768, n_8769, n_8770, n_8771, n_8772, n_8773, n_8774,
          n_8775, n_8776, a_SMASKREG_F2_G_aNOT_aCLK, a_N2571_aNOT, a_EQ624,
          n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, a_SCOMMANDREG_F2_G,
          a_SCOMMANDREG_F2_G_aCLRN, a_EQ1125, n_8793, n_8794, n_8795, n_8796,
          n_8797, n_8798, n_8799, n_8800, n_8801, n_8802, a_SCOMMANDREG_F2_G_aCLK,
          a_LC5_B8_aNOT, a_EQ466, n_8806, n_8807, n_8808, n_8809, n_8810,
          n_8811, n_8812, a_N1565, a_EQ464, n_8815, n_8816, n_8817, n_8818,
          n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, a_LC4_B8, a_EQ467,
          n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833, n_8834,
          n_8835, a_N1563_aNOT, a_EQ463, n_8838, n_8839, n_8840, n_8841, a_SMASKREG_F3_G_aNOT,
          n_8843, n_8844, n_8845, n_8846, n_8847, a_N24, a_EQ177, n_8850,
          n_8851, n_8852, n_8853, n_8854, n_8855, n_8856, n_8857, a_LC2_B8_aNOT,
          a_EQ461, n_8860, n_8861, n_8862, n_8863, n_8864, n_8865, n_8866,
          n_8867, a_LC1_B8, a_EQ462, n_8870, n_8871, n_8872, n_8873, n_8874,
          n_8875, n_8876, n_8877, n_8878, a_SMASKREG_F3_G_aNOT_aCLRN, a_EQ1160,
          n_8885, n_8886, n_8887, n_8888, n_8889, n_8890, n_8891, n_8892,
          n_8893, n_8894, a_SMASKREG_F3_G_aNOT_aCLK, a_STCSTATUS_F3_G, a_STCSTATUS_F3_G_aCLRN,
          a_EQ1180, n_8903, n_8904, n_8905, n_8906, n_8907, n_8908, n_8909,
          n_8910, n_8911, n_8912, a_STCSTATUS_F3_G_aCLK, a_LC3_B18, a_EQ541,
          n_8916, n_8917, n_8918, a_SREQUESTREG_F3_G, n_8920, n_8921, n_8922,
          n_8923, n_8924, a_SREQUESTREG_F3_G_aCLRN, a_EQ1176, n_8931, n_8932,
          n_8933, n_8934, n_8935, n_8936, n_8937, n_8938, n_8939, n_8940,
          n_8941, a_SREQUESTREG_F3_G_aCLK, a_SCOMMANDREG_F3_G, a_SCOMMANDREG_F3_G_aCLRN,
          a_EQ1126, n_8950, n_8951, n_8952, n_8953, n_8954, n_8955, n_8956,
          n_8957, n_8958, n_8959, a_SCOMMANDREG_F3_G_aCLK, a_SCOMMANDREG_F4_G,
          a_SCOMMANDREG_F4_G_aCLRN, a_EQ1127, n_8968, n_8969, n_8970, n_8971,
          n_8972, n_8973, n_8974, n_8975, n_8976, n_8977, a_SCOMMANDREG_F4_G_aCLK,
          a_SCH3MODEREG_F5_G, a_SCH3MODEREG_F5_G_aCLRN, a_EQ1112, n_8986,
          n_8987, n_8988, n_8989, n_8990, n_8991, n_8992, n_8993, n_8994,
          a_SCH3MODEREG_F5_G_aCLK, a_SCH1MODEREG_F5_G, a_SCH1MODEREG_F5_G_aCLRN,
          a_EQ984, n_9003, n_9004, n_9005, n_9006, n_9007, n_9008, n_9009,
          n_9010, n_9011, a_SCH1MODEREG_F5_G_aCLK, a_SCH2MODEREG_F5_G, a_SCH2MODEREG_F5_G_aCLRN,
          a_EQ1048, n_9020, n_9021, n_9022, n_9023, n_9024, n_9025, n_9026,
          n_9027, n_9028, a_SCH2MODEREG_F5_G_aCLK, a_LC1_B15, a_EQ533, n_9032,
          n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040,
          n_9041, n_9042, a_N2390, a_N2390_aIN, n_9045, n_9046, n_9047, n_9048,
          n_9049, a_SMODECOUNTER_F1_G, a_SMODECOUNTER_F1_G_aCLRN, a_EQ1162,
          n_9057, n_9058, n_9059, n_9060, n_9061, a_SMODECOUNTER_F0_G, n_9063,
          n_9064, n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071,
          n_9072, n_9073, a_SMODECOUNTER_F1_G_aCLK, a_SMODECOUNTER_F0_G_aCLRN,
          a_EQ1161, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087,
          n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095,
          n_9096, a_SMODECOUNTER_F0_G_aCLK, a_SCH0MODEREG_F5_G, a_SCH0MODEREG_F5_G_aCLRN,
          a_EQ920, n_9105, n_9106, n_9107, n_9108, n_9109, n_9110, n_9111,
          n_9112, n_9113, a_SCH0MODEREG_F5_G_aCLK, a_SCH2BAROUT_F0_G, a_SCH2BAROUT_F0_G_aCLRN,
          a_EQ1011, n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128,
          n_9129, n_9130, a_SCH2BAROUT_F0_G_aCLK, a_SCH2MODEREG_F2_G_aCLRN,
          a_EQ1045, n_9138, n_9139, n_9140, n_9141, n_9142, n_9143, n_9144,
          n_9145, n_9146, a_SCH2MODEREG_F2_G_aCLK, a_SCH3BAROUT_F0_G, a_SCH3BAROUT_F0_G_aCLRN,
          a_EQ1075, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160, n_9161,
          n_9162, n_9163, a_SCH3BAROUT_F0_G_aCLK, a_SCH3MODEREG_F2_G_aCLRN,
          a_EQ1109, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176, n_9177,
          n_9178, n_9179, a_SCH3MODEREG_F2_G_aCLK, a_SCH0BAROUT_F0_G, a_SCH0BAROUT_F0_G_aCLRN,
          a_EQ883, n_9188, n_9189, n_9190, n_9191, n_9192, n_9193, n_9194,
          n_9195, n_9196, a_SCH0BAROUT_F0_G_aCLK, a_N2584_aNOT, a_EQ637, n_9200,
          n_9201, n_9202, n_9203, n_9204, n_9205, a_SCH1BAROUT_F0_G, a_SCH1BAROUT_F0_G_aCLRN,
          a_EQ947, n_9213, n_9214, n_9215, n_9216, n_9217, n_9218, n_9219,
          n_9220, n_9221, a_SCH1BAROUT_F0_G_aCLK, a_SCOMMANDREG_F1_G_aCLRN,
          a_EQ1124, n_9229, n_9230, n_9231, n_9232, n_9233, n_9234, n_9235,
          n_9236, n_9237, n_9238, a_SCOMMANDREG_F1_G_aCLK, a_SCH1BAROUT_F1_G,
          a_SCH1BAROUT_F1_G_aCLRN, a_EQ948, n_9247, n_9248, n_9249, n_9250,
          n_9251, n_9252, n_9253, n_9254, n_9255, a_SCH1BAROUT_F1_G_aCLK,
          a_SCH0BAROUT_F1_G, a_SCH0BAROUT_F1_G_aCLRN, a_EQ884, n_9264, n_9265,
          n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, a_SCH0BAROUT_F1_G_aCLK,
          a_SCH3BAROUT_F1_G, a_SCH3BAROUT_F1_G_aCLRN, a_EQ1076, n_9281, n_9282,
          n_9283, n_9284, n_9285, n_9286, n_9287, n_9288, n_9289, a_SCH3BAROUT_F1_G_aCLK,
          a_SCH1BAROUT_F2_G, a_SCH1BAROUT_F2_G_aCLRN, a_EQ949, n_9298, n_9299,
          n_9300, n_9301, n_9302, n_9303, n_9304, n_9305, n_9306, a_SCH1BAROUT_F2_G_aCLK,
          a_SCH3BAROUT_F2_G, a_SCH3BAROUT_F2_G_aCLRN, a_EQ1077, n_9315, n_9316,
          n_9317, n_9318, n_9319, n_9320, n_9321, n_9322, n_9323, a_SCH3BAROUT_F2_G_aCLK,
          a_SCH2BAROUT_F2_G, a_SCH2BAROUT_F2_G_aCLRN, a_EQ1013, n_9332, n_9333,
          n_9334, n_9335, n_9336, n_9337, n_9338, n_9339, n_9340, a_SCH2BAROUT_F2_G_aCLK,
          a_SCH0BAROUT_F2_G, a_SCH0BAROUT_F2_G_aCLRN, a_EQ885, n_9349, n_9350,
          n_9351, n_9352, n_9353, n_9354, n_9355, n_9356, n_9357, a_SCH0BAROUT_F2_G_aCLK,
          a_SCH0BAROUT_F3_G, a_SCH0BAROUT_F3_G_aCLRN, a_EQ886, n_9366, n_9367,
          n_9368, n_9369, n_9370, n_9371, n_9372, n_9373, n_9374, a_SCH0BAROUT_F3_G_aCLK,
          a_SCH2BAROUT_F3_G, a_SCH2BAROUT_F3_G_aCLRN, a_EQ1014, n_9383, n_9384,
          n_9385, n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, a_SCH2BAROUT_F3_G_aCLK,
          a_SCH1BAROUT_F3_G, a_SCH1BAROUT_F3_G_aCLRN, a_EQ950, n_9400, n_9401,
          n_9402, n_9403, n_9404, n_9405, n_9406, n_9407, n_9408, a_SCH1BAROUT_F3_G_aCLK,
          a_SCH3BAROUT_F3_G, a_SCH3BAROUT_F3_G_aCLRN, a_EQ1078, n_9417, n_9418,
          n_9419, n_9420, n_9421, n_9422, n_9423, n_9424, n_9425, a_SCH3BAROUT_F3_G_aCLK,
          a_SCH1BAROUT_F4_G, a_SCH1BAROUT_F4_G_aCLRN, a_EQ951, n_9434, n_9435,
          n_9436, n_9437, n_9438, n_9439, n_9440, n_9441, n_9442, a_SCH1BAROUT_F4_G_aCLK,
          a_SCH2BAROUT_F4_G, a_SCH2BAROUT_F4_G_aCLRN, a_EQ1015, n_9451, n_9452,
          n_9453, n_9454, n_9455, n_9456, n_9457, n_9458, n_9459, a_SCH2BAROUT_F4_G_aCLK,
          a_SCH3BAROUT_F4_G, a_SCH3BAROUT_F4_G_aCLRN, a_EQ1079, n_9468, n_9469,
          n_9470, n_9471, n_9472, n_9473, n_9474, n_9475, n_9476, a_SCH3BAROUT_F4_G_aCLK,
          a_SCH0BAROUT_F4_G, a_SCH0BAROUT_F4_G_aCLRN, a_EQ887, n_9485, n_9486,
          n_9487, n_9488, n_9489, n_9490, n_9491, n_9492, n_9493, a_SCH0BAROUT_F4_G_aCLK,
          a_SCH1BAROUT_F5_G, a_SCH1BAROUT_F5_G_aCLRN, a_EQ952, n_9502, n_9503,
          n_9504, n_9505, n_9506, n_9507, n_9508, n_9509, n_9510, a_SCH1BAROUT_F5_G_aCLK,
          a_SCH2BAROUT_F5_G, a_SCH2BAROUT_F5_G_aCLRN, a_EQ1016, n_9519, n_9520,
          n_9521, n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, a_SCH2BAROUT_F5_G_aCLK,
          a_SCH0BAROUT_F5_G, a_SCH0BAROUT_F5_G_aCLRN, a_EQ888, n_9536, n_9537,
          n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, a_SCH0BAROUT_F5_G_aCLK,
          a_SCH2BAROUT_F6_G, a_SCH2BAROUT_F6_G_aCLRN, a_EQ1017, n_9553, n_9554,
          n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561, a_SCH2BAROUT_F6_G_aCLK,
          a_SCH0BAROUT_F6_G, a_SCH0BAROUT_F6_G_aCLRN, a_EQ889, n_9570, n_9571,
          n_9572, n_9573, n_9574, n_9575, n_9576, n_9577, n_9578, a_SCH0BAROUT_F6_G_aCLK,
          a_SCH1BAROUT_F6_G, a_SCH1BAROUT_F6_G_aCLRN, a_EQ953, n_9587, n_9588,
          n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, a_SCH1BAROUT_F6_G_aCLK,
          a_SCH3BAROUT_F6_G, a_SCH3BAROUT_F6_G_aCLRN, a_EQ1081, n_9604, n_9605,
          n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612, a_SCH3BAROUT_F6_G_aCLK,
          a_SCH2BAROUT_F7_G, a_SCH2BAROUT_F7_G_aCLRN, a_EQ1018, n_9621, n_9622,
          n_9623, n_9624, n_9625, n_9626, n_9627, n_9628, n_9629, a_SCH2BAROUT_F7_G_aCLK,
          a_SCH0MODEREG_F2_G_aCLRN, a_EQ917, n_9637, n_9638, n_9639, n_9640,
          n_9641, n_9642, n_9643, n_9644, n_9645, a_SCH0MODEREG_F2_G_aCLK,
          a_SCH0BAROUT_F7_G, a_SCH0BAROUT_F7_G_aCLRN, a_EQ890, n_9654, n_9655,
          n_9656, n_9657, n_9658, n_9659, n_9660, n_9661, n_9662, a_SCH0BAROUT_F7_G_aCLK,
          a_SCH1MODEREG_F2_G_aCLRN, a_EQ981, n_9670, n_9671, n_9672, n_9673,
          n_9674, n_9675, n_9676, n_9677, n_9678, a_SCH1MODEREG_F2_G_aCLK,
          a_SCH1BAROUT_F7_G, a_SCH1BAROUT_F7_G_aCLRN, a_EQ954, n_9687, n_9688,
          n_9689, n_9690, n_9691, n_9692, n_9693, n_9694, n_9695, a_SCH1BAROUT_F7_G_aCLK,
          a_SCH2MODEREG_F0_G_aCLRN, a_EQ1043, n_9703, n_9704, n_9705, n_9706,
          n_9707, n_9708, n_9709, n_9710, n_9711, a_SCH2MODEREG_F0_G_aCLK,
          a_SCH1MODEREG_F0_G_aCLRN, a_EQ979, n_9719, n_9720, n_9721, n_9722,
          n_9723, n_9724, n_9725, n_9726, n_9727, a_SCH1MODEREG_F0_G_aCLK,
          a_SCH0MODEREG_F0_G_aCLRN, a_EQ915, n_9735, n_9736, n_9737, n_9738,
          n_9739, n_9740, n_9741, n_9742, n_9743, a_SCH0MODEREG_F0_G_aCLK,
          a_SCH3MODEREG_F0_G_aCLRN, a_EQ1107, n_9751, n_9752, n_9753, n_9754,
          n_9755, n_9756, n_9757, n_9758, n_9759, a_SCH3MODEREG_F0_G_aCLK,
          a_SCH1MODEREG_F1_G_aCLRN, a_EQ980, n_9767, n_9768, n_9769, n_9770,
          n_9771, n_9772, n_9773, n_9774, n_9775, a_SCH1MODEREG_F1_G_aCLK,
          a_SCH3MODEREG_F1_G_aCLRN, a_EQ1108, n_9783, n_9784, n_9785, n_9786,
          n_9787, n_9788, n_9789, n_9790, n_9791, a_SCH3MODEREG_F1_G_aCLK,
          a_SCH0MODEREG_F1_G_aCLRN, a_EQ916, n_9799, n_9800, n_9801, n_9802,
          n_9803, n_9804, n_9805, n_9806, n_9807, a_SCH0MODEREG_F1_G_aCLK,
          a_SCH2MODEREG_F1_G_aCLRN, a_EQ1044, n_9815, n_9816, n_9817, n_9818,
          n_9819, n_9820, n_9821, n_9822, n_9823, a_SCH2MODEREG_F1_G_aCLK,
          a_LC2_E21, a_EQ375, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832,
          n_9833, n_9834, a_N1162_aNOT, a_EQ372, n_9837, n_9838, n_9839, n_9840,
          n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848,
          a_N1168, a_EQ377, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856,
          n_9857, n_9858, a_N1169, a_EQ378, n_9861, n_9862, n_9863, n_9864,
          n_9865, n_9866, n_9867, n_9868, n_9869, n_9870, a_LC3_E21, a_EQ376,
          n_9873, n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880,
          a_N3546_aCLRN, a_EQ842, n_9887, n_9888, n_9889, n_9890, n_9891,
          n_9892, n_9893, n_9894, n_9895, n_9896, n_9897, n_9898, a_N3546_aCLK,
          a_LC4_A20, a_EQ259, n_9902, n_9903, n_9904, n_9905, n_9906, n_9907,
          n_9908, n_9909, n_9910, n_9911, n_9912, n_9913, n_9914, n_9915,
          n_9916, n_9917, a_LC2_A20, a_EQ258, n_9920, n_9921, n_9922, n_9923,
          n_9924, n_9925, n_9926, n_9927, a_N517_aNOT, a_EQ262, n_9930, n_9931,
          n_9932, n_9933, n_9934, n_9935, n_9936, n_9937, a_LC8_A26, a_EQ261,
          n_9940, n_9941, n_9942, n_9943, n_9944, n_9945, n_9946, n_9947,
          a_LC8_A20, a_EQ260, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955,
          n_9956, n_9957, a_N3545_aCLRN, a_EQ841, n_9964, n_9965, n_9966,
          n_9967, n_9968, n_9969, n_9970, n_9971, n_9972, n_9973, n_9974,
          n_9975, a_N3545_aCLK, a_LC3_A1, a_EQ403, n_9979, n_9980, n_9981,
          n_9982, n_9983, n_9984, n_9985, n_9986, a_N1297_aNOT, a_EQ410, n_9989,
          n_9990, n_9991, n_9992, n_9993, n_9994, n_9995, n_9996, a_N1286,
          a_EQ402, n_9999, n_10000, n_10001, n_10002, n_10003, n_10004, n_10005,
          n_10006, a_N1285, a_EQ401, n_10009, n_10010, n_10011, n_10012, n_10013,
          n_10014, n_10015, n_10016, n_10017, n_10018, a_LC1_A1, a_EQ404,
          n_10021, n_10022, n_10023, n_10024, n_10025, n_10026, n_10027, n_10028,
          a_N3544_aCLRN, a_EQ840, n_10035, n_10036, n_10037, n_10038, n_10039,
          n_10040, n_10041, n_10042, n_10043, n_10044, n_10045, n_10046, a_N3544_aCLK,
          a_LC7_E14, a_EQ340, n_10051, n_10052, n_10053, n_10054, n_10055,
          n_10056, n_10057, n_10058, a_LC4_E14, a_EQ339, n_10061, n_10062,
          n_10063, n_10064, n_10065, n_10066, n_10067, n_10068, a_N1019_aNOT,
          a_EQ341, n_10071, n_10072, n_10073, n_10074, n_10075, n_10076, n_10077,
          n_10078, a_LC5_E14, a_EQ338, n_10081, n_10082, n_10083, n_10084,
          n_10085, n_10086, n_10087, n_10088, a_LC6_E14, a_EQ337, n_10091,
          n_10092, n_10093, n_10094, n_10095, n_10096, n_10097, n_10098, a_SADDRESSOUT_F13_G_aCLRN,
          a_EQ859, n_10105, n_10106, n_10107, n_10108, n_10109, n_10110, n_10111,
          n_10112, n_10113, n_10114, n_10115, n_10116, a_SADDRESSOUT_F13_G_aCLK,
          a_LC7_D6, a_EQ407, n_10120, n_10121, n_10122, n_10123, n_10124,
          n_10125, n_10126, n_10127, a_N1298_aNOT, a_EQ411, n_10130, n_10131,
          n_10132, n_10133, n_10134, n_10135, n_10136, n_10137, a_N1292, a_EQ406,
          n_10140, n_10141, n_10142, n_10143, n_10144, n_10145, n_10146, n_10147,
          a_N1291, a_EQ405, n_10150, n_10151, n_10152, n_10153, n_10154, n_10155,
          n_10156, n_10157, n_10158, n_10159, a_LC1_D14, a_EQ408, n_10162,
          n_10163, n_10164, n_10165, n_10166, n_10167, n_10168, n_10169, a_SADDRESSOUT_F15_G_aCLRN,
          a_EQ861, n_10176, n_10177, n_10178, n_10179, n_10180, n_10181, n_10182,
          n_10183, n_10184, n_10185, n_10186, n_10187, a_SADDRESSOUT_F15_G_aCLK,
          a_EQ1132, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195,
          n_10196, n_10197, a_N825_aCLRN, a_EQ310, n_10205, n_10206, n_10207,
          n_10208, n_10209, n_10210, n_10211, n_10212, n_10213, a_N825_aCLK,
          a_LC6_E3, a_EQ233, n_10217, n_10218, n_10219, n_10220, n_10221,
          n_10222, n_10223, n_10224, n_10225, n_10226, n_10227, n_10228, a_LC4_E3,
          a_EQ232, n_10231, n_10232, n_10233, n_10234, n_10235, n_10236, n_10237,
          n_10238, a_N340_aNOT, a_EQ234, n_10241, n_10242, n_10243, n_10244,
          n_10245, n_10246, n_10247, n_10248, a_LC3_E3, a_EQ231, n_10251,
          n_10252, n_10253, n_10254, n_10255, n_10256, n_10257, n_10258, a_LC2_E3,
          a_EQ230, n_10261, n_10262, n_10263, n_10264, n_10265, n_10266, n_10267,
          n_10268, a_N3543_aCLRN, a_EQ839, n_10275, n_10276, n_10277, n_10278,
          n_10279, n_10280, n_10281, n_10282, n_10283, n_10284, n_10285, n_10286,
          a_N3543_aCLK, a_N866_aNOT, a_EQ317, n_10290, n_10291, n_10292, n_10293,
          n_10294, n_10295, n_10296, n_10297, n_10298, n_10299, n_10300, n_10301,
          n_10302, n_10303, n_10304, n_10305, a_N874, a_EQ321, n_10308, n_10309,
          n_10310, n_10311, n_10312, n_10313, n_10314, n_10315, a_LC8_E16,
          a_EQ322, n_10318, n_10319, n_10320, n_10321, n_10322, n_10323, n_10324,
          n_10325, a_LC2_E16, a_EQ320, n_10328, n_10329, n_10330, n_10331,
          n_10332, n_10333, n_10334, n_10335, a_LC1_E16, a_EQ319, n_10338,
          n_10339, n_10340, n_10341, n_10342, n_10343, n_10344, n_10345, a_N3542_aCLRN,
          a_EQ838, n_10352, n_10353, n_10354, n_10355, n_10356, n_10357, n_10358,
          n_10359, n_10360, n_10361, n_10362, n_10363, a_N3542_aCLK, a_N2372_aNOT,
          a_N2372_aNOT_aIN, n_10367, n_10368, n_10369, n_10370, n_10371, n_10372,
          n_10373, a_STEMPORARYREG_F0_G, a_STEMPORARYREG_F0_G_aCLRN, a_EQ1181,
          n_10381, n_10382, n_10383, n_10384, n_10385, n_10386, n_10387, n_10388,
          n_10389, n_10390, n_10391, a_STEMPORARYREG_F0_G_aCLK, a_N1338_aNOT,
          a_EQ425, n_10395, n_10396, n_10397, n_10398, n_10399, n_10400, n_10401,
          n_10402, a_N1327, a_EQ417, n_10405, n_10406, n_10407, n_10408, n_10409,
          n_10410, n_10411, n_10412, a_LC6_F5, a_EQ416, n_10415, n_10416,
          n_10417, n_10418, n_10419, n_10420, n_10421, n_10422, a_LC1_F5,
          a_EQ419, n_10425, n_10426, n_10427, n_10428, n_10429, n_10430, n_10431,
          n_10432, a_LC2_F5, a_EQ418, n_10435, n_10436, n_10437, n_10438,
          n_10439, n_10440, n_10441, n_10442, a_SADDRESSOUT_F8_G_aCLRN, a_EQ854,
          n_10449, n_10450, n_10451, n_10452, n_10453, n_10454, n_10455, n_10456,
          n_10457, n_10458, n_10459, n_10460, a_SADDRESSOUT_F8_G_aCLK, a_SCOMMANDREG_F0_G_aCLRN,
          a_EQ1123, n_10468, n_10469, n_10470, n_10471, n_10472, n_10473,
          n_10474, n_10475, n_10476, n_10477, n_10478, a_SCOMMANDREG_F0_G_aCLK,
          a_STEMPORARYREG_F1_G, a_STEMPORARYREG_F1_G_aCLRN, a_EQ1182, n_10487,
          n_10488, n_10489, n_10490, n_10491, n_10492, n_10493, n_10494, n_10495,
          n_10496, n_10497, a_STEMPORARYREG_F1_G_aCLK, a_LC2_A18, a_EQ279,
          n_10501, n_10502, n_10503, n_10504, n_10505, n_10506, n_10507, n_10508,
          a_LC1_A18, a_EQ280, n_10511, n_10512, n_10513, n_10514, n_10515,
          n_10516, n_10517, n_10518, a_N672_aNOT, a_EQ283, n_10521, n_10522,
          n_10523, n_10524, n_10525, n_10526, n_10527, n_10528, a_LC4_A18,
          a_EQ282, n_10531, n_10532, n_10533, n_10534, n_10535, n_10536, n_10537,
          n_10538, a_LC5_A18, a_EQ281, n_10541, n_10542, n_10543, n_10544,
          n_10545, n_10546, n_10547, n_10548, a_SADDRESSOUT_F9_G_aCLRN, a_EQ855,
          n_10555, n_10556, n_10557, n_10558, n_10559, n_10560, n_10561, n_10562,
          n_10563, n_10564, n_10565, n_10566, a_SADDRESSOUT_F9_G_aCLK, a_LC3_E15,
          a_EQ333, n_10570, n_10571, n_10572, n_10573, n_10574, n_10575, n_10576,
          n_10577, a_LC1_E18, a_EQ332, n_10580, n_10581, n_10582, n_10583,
          n_10584, n_10585, n_10586, n_10587, a_N1000_aNOT, a_EQ336, n_10590,
          n_10591, n_10592, n_10593, n_10594, n_10595, n_10596, n_10597, a_LC1_E21,
          a_EQ335, n_10600, n_10601, n_10602, n_10603, n_10604, n_10605, n_10606,
          n_10607, a_LC8_E15, a_EQ334, n_10610, n_10611, n_10612, n_10613,
          n_10614, n_10615, n_10616, n_10617, a_SADDRESSOUT_F10_G_aCLRN, a_EQ856,
          n_10624, n_10625, n_10626, n_10627, n_10628, n_10629, n_10630, n_10631,
          n_10632, n_10633, n_10634, n_10635, a_SADDRESSOUT_F10_G_aCLK, a_STEMPORARYREG_F2_G,
          a_STEMPORARYREG_F2_G_aCLRN, a_EQ1183, n_10644, n_10645, n_10646,
          n_10647, n_10648, n_10649, n_10650, n_10651, n_10652, n_10653, n_10654,
          a_STEMPORARYREG_F2_G_aCLK, a_N1339_aNOT, a_EQ426, n_10658, n_10659,
          n_10660, n_10661, n_10662, n_10663, n_10664, n_10665, a_N1333, a_EQ421,
          n_10668, n_10669, n_10670, n_10671, n_10672, n_10673, n_10674, n_10675,
          a_LC3_A19, a_EQ420, n_10678, n_10679, n_10680, n_10681, n_10682,
          n_10683, n_10684, n_10685, a_LC1_A19, a_EQ423, n_10688, n_10689,
          n_10690, n_10691, n_10692, n_10693, n_10694, n_10695, a_LC2_A19,
          a_EQ422, n_10698, n_10699, n_10700, n_10701, n_10702, n_10703, n_10704,
          n_10705, a_SADDRESSOUT_F11_G_aCLRN, a_EQ857, n_10712, n_10713, n_10714,
          n_10715, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721, n_10722,
          n_10723, a_SADDRESSOUT_F11_G_aCLK, a_STEMPORARYREG_F3_G, a_STEMPORARYREG_F3_G_aCLRN,
          a_EQ1184, n_10732, n_10733, n_10734, n_10735, n_10736, n_10737,
          n_10738, n_10739, n_10740, n_10741, n_10742, a_STEMPORARYREG_F3_G_aCLK,
          a_LC3_A26, a_EQ207, n_10746, n_10747, n_10748, n_10749, n_10750,
          n_10751, n_10752, n_10753, a_LC2_A26, a_EQ206, n_10756, n_10757,
          n_10758, n_10759, n_10760, n_10761, n_10762, n_10763, a_LC4_A26,
          a_EQ210, n_10766, n_10767, n_10768, n_10769, n_10770, n_10771, n_10772,
          n_10773, a_LC5_A26, a_EQ209, n_10776, n_10777, n_10778, n_10779,
          n_10780, n_10781, n_10782, n_10783, a_LC6_A26, a_EQ208, n_10786,
          n_10787, n_10788, n_10789, n_10790, n_10791, n_10792, n_10793, a_SADDRESSOUT_F12_G_aCLRN,
          a_EQ858, n_10800, n_10801, n_10802, n_10803, n_10804, n_10805, n_10806,
          n_10807, n_10808, n_10809, n_10810, n_10811, a_SADDRESSOUT_F12_G_aCLK,
          a_SCOMMANDREG_F6_G, a_SCOMMANDREG_F6_G_aCLRN, a_EQ1129, n_10820,
          n_10821, n_10822, n_10823, n_10824, n_10825, n_10826, n_10827, n_10828,
          n_10829, a_SCOMMANDREG_F6_G_aCLK, a_STEMPORARYREG_F5_G, a_STEMPORARYREG_F5_G_aCLRN,
          a_EQ1186, n_10838, n_10839, n_10840, n_10841, n_10842, n_10843,
          n_10844, n_10845, n_10846, n_10847, n_10848, a_STEMPORARYREG_F5_G_aCLK,
          a_STEMPORARYREG_F6_G, a_STEMPORARYREG_F6_G_aCLRN, a_EQ1187, n_10857,
          n_10858, n_10859, n_10860, n_10861, n_10862, n_10863, n_10864, n_10865,
          n_10866, n_10867, a_STEMPORARYREG_F6_G_aCLK, a_LC4_F9, a_EQ218,
          n_10871, n_10872, n_10873, n_10874, n_10875, n_10876, n_10877, n_10878,
          a_LC7_F9, a_EQ217, n_10881, n_10882, n_10883, n_10884, n_10885,
          n_10886, n_10887, n_10888, a_N240_aNOT, a_EQ219, n_10891, n_10892,
          n_10893, n_10894, n_10895, n_10896, n_10897, n_10898, a_LC3_F9,
          a_EQ216, n_10901, n_10902, n_10903, n_10904, n_10905, n_10906, n_10907,
          n_10908, a_LC1_F9, a_EQ215, n_10911, n_10912, n_10913, n_10914,
          n_10915, n_10916, n_10917, n_10918, a_SADDRESSOUT_F14_G_aCLRN, a_EQ860,
          n_10925, n_10926, n_10927, n_10928, n_10929, n_10930, n_10931, n_10932,
          n_10933, n_10934, n_10935, n_10936, a_SADDRESSOUT_F14_G_aCLK, a_N1776_aNOT,
          a_EQ508, n_10940, n_10941, n_10942, n_10943, n_10944, n_10945, n_10946,
          n_10947, a_LC6_A4, a_LC6_A4_aIN, n_10950, n_10951, n_10952, n_10953,
          n_10954, n_10955, bytepointer_aCLRN, a_EQ001, n_10962, n_10963,
          n_10964, n_10965, n_10966, n_10967, n_10968, n_10969, n_10970, bytepointer_aCLK,
          a_STEMPORARYREG_F7_G, a_STEMPORARYREG_F7_G_aCLRN, a_EQ1188, n_10979,
          n_10980, n_10981, n_10982, n_10983, n_10984, n_10985, n_10986, n_10987,
          n_10988, n_10989, a_STEMPORARYREG_F7_G_aCLK, a_LC2_F19, a_EQ285,
          n_10993, n_10994, n_10995, n_10996, a_SCH2ADDRREG_F0_G, n_10998,
          n_10999, n_11000, n_11001, n_11002, n_11003, n_11004, n_11005, a_LC3_F19,
          a_EQ723, n_11008, n_11009, n_11010, n_11011, n_11012, n_11013, n_11014,
          n_11015, n_11016, n_11017, n_11018, n_11019, a_SCH2ADDRREG_F0_G_aCLRN,
          a_EQ995, n_11026, n_11027, n_11028, n_11029, n_11030, n_11031, n_11032,
          n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, a_SCH2ADDRREG_F0_G_aCLK,
          a_N1493_aNOT, a_EQ455, n_11042, n_11043, n_11044, n_11045, a_SCH3ADDRREG_F0_G,
          n_11047, n_11048, n_11049, n_11050, n_11051, n_11052, n_11053, n_11054,
          a_LC8_D8, a_EQ456, n_11057, n_11058, n_11059, n_11060, n_11061,
          n_11062, n_11063, n_11064, n_11065, n_11066, n_11067, n_11068, a_SCH3ADDRREG_F0_G_aCLRN,
          a_EQ1059, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080,
          n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087, a_SCH3ADDRREG_F0_G_aCLK,
          a_LC1_D8, a_EQ673, n_11091, n_11092, n_11093, n_11094, a_SCH0ADDRREG_F0_G,
          n_11096, n_11097, n_11098, n_11099, n_11100, n_11101, n_11102, n_11103,
          a_LC4_D8, a_EQ674, n_11106, n_11107, n_11108, n_11109, n_11110,
          n_11111, n_11112, n_11113, n_11114, n_11115, n_11116, n_11117, n_11118,
          a_SCH0ADDRREG_F0_G_aCLRN, a_EQ867, n_11125, n_11126, n_11127, n_11128,
          n_11129, n_11130, n_11131, n_11132, n_11133, n_11134, n_11135, n_11136,
          n_11137, a_SCH0ADDRREG_F0_G_aCLK, a_LC2_D19, a_EQ698, n_11141, n_11142,
          n_11143, n_11144, a_SCH1ADDRREG_F0_G, n_11146, n_11147, n_11148,
          n_11149, n_11150, n_11151, n_11152, n_11153, a_LC1_D19, a_EQ699,
          n_11156, n_11157, n_11158, n_11159, n_11160, n_11161, n_11162, n_11163,
          n_11164, n_11165, n_11166, n_11167, n_11168, a_SCH1ADDRREG_F0_G_aCLRN,
          a_EQ931, n_11175, n_11176, n_11177, n_11178, n_11179, n_11180, n_11181,
          n_11182, n_11183, n_11184, n_11185, n_11186, n_11187, a_SCH1ADDRREG_F0_G_aCLK,
          a_N3059, a_EQ836, n_11191, n_11192, n_11193, n_11194, n_11195, n_11196,
          n_11197, n_11198, n_11199, n_11200, n_11201, n_11202, n_11203, n_11204,
          n_11205, n_11206, n_11207, n_11208, a_LC3_C9, a_EQ235, n_11211,
          n_11212, n_11213, n_11214, n_11215, n_11216, n_11217, n_11218, n_11219,
          n_11220, a_LC2_C9, a_EQ697, n_11223, n_11224, n_11225, n_11226,
          n_11227, n_11228, n_11229, n_11230, n_11231, a_SCH1ADDRREG_F1_G,
          n_11233, a_SCH1ADDRREG_F1_G_aCLRN, a_EQ932, n_11240, n_11241, n_11242,
          n_11243, n_11244, n_11245, n_11246, n_11247, n_11248, n_11249, n_11250,
          n_11251, a_SCH1ADDRREG_F1_G_aCLK, a_LC4_C9, a_EQ270, n_11255, n_11256,
          n_11257, n_11258, n_11259, n_11260, n_11261, n_11262, n_11263, n_11264,
          a_LC5_C9, a_EQ672, n_11267, n_11268, n_11269, n_11270, n_11271,
          n_11272, n_11273, n_11274, n_11275, a_SCH0ADDRREG_F1_G, n_11277,
          a_SCH0ADDRREG_F1_G_aCLRN, a_EQ868, n_11284, n_11285, n_11286, n_11287,
          n_11288, n_11289, n_11290, n_11291, n_11292, n_11293, n_11294, n_11295,
          a_SCH0ADDRREG_F1_G_aCLK, a_LC3_C12, a_EQ721, n_11299, n_11300, n_11301,
          n_11302, n_11303, n_11304, n_11305, n_11306, n_11307, a_LC5_C12,
          a_EQ722, n_11310, n_11311, n_11312, n_11313, n_11314, n_11315, n_11316,
          n_11317, a_SCH2ADDRREG_F1_G, a_SCH2ADDRREG_F1_G_aCLRN, a_EQ996,
          n_11325, n_11326, n_11327, n_11328, n_11329, n_11330, n_11331, n_11332,
          n_11333, a_SCH2ADDRREG_F1_G_aCLK, a_N937_aNOT, a_N937_aNOT_aIN,
          n_11337, n_11338, n_11339, n_11340, n_11341, a_LC2_C26, a_EQ747,
          n_11344, n_11345, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351,
          n_11352, a_SCH3ADDRREG_F1_G, n_11354, a_SCH3ADDRREG_F1_G_aCLRN,
          a_EQ1060, n_11361, n_11362, n_11363, n_11364, n_11365, n_11366,
          n_11367, n_11368, n_11369, n_11370, a_SCH3ADDRREG_F1_G_aCLK, a_N2542,
          a_EQ599, n_11374, n_11375, n_11376, n_11377, n_11378, n_11379, n_11380,
          n_11381, n_11382, n_11383, n_11384, n_11385, n_11386, a_LC1_C2,
          a_EQ695, n_11389, n_11390, n_11391, n_11392, a_SCH1ADDRREG_F2_G,
          n_11394, n_11395, n_11396, n_11397, n_11398, n_11399, n_11400, n_11401,
          a_LC2_C2, a_EQ696, n_11404, n_11405, n_11406, n_11407, n_11408,
          n_11409, n_11410, n_11411, a_SCH1ADDRREG_F2_G_aCLRN, a_EQ933, n_11418,
          n_11419, n_11420, n_11421, n_11422, n_11423, n_11424, n_11425, n_11426,
          n_11427, n_11428, n_11429, n_11430, a_SCH1ADDRREG_F2_G_aCLK, a_N930_aNOT,
          a_EQ325, n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440,
          n_11441, n_11442, n_11443, a_LC5_C20, a_EQ746, n_11446, n_11447,
          n_11448, n_11449, n_11450, n_11451, n_11452, n_11453, n_11454, a_SCH3ADDRREG_F2_G,
          n_11456, a_SCH3ADDRREG_F2_G_aCLRN, a_EQ1061, n_11463, n_11464, n_11465,
          n_11466, n_11467, n_11468, n_11469, n_11470, n_11471, n_11472, a_SCH3ADDRREG_F2_G_aCLK,
          a_N740_aNOT, a_N740_aNOT_aIN, n_11476, n_11477, n_11478, n_11479,
          n_11480, n_11481, a_SCH2ADDRREG_F2_G, n_11483, a_N2434, a_N2434_aIN,
          n_11486, n_11487, n_11488, n_11489, n_11490, a_LC4_C5, a_EQ720,
          n_11493, n_11494, n_11495, n_11496, n_11497, n_11498, n_11499, n_11500,
          n_11501, n_11502, n_11503, n_11504, n_11505, a_SCH2ADDRREG_F2_G_aCLRN,
          a_EQ997, n_11512, n_11513, n_11514, n_11515, n_11516, n_11517, n_11518,
          n_11519, n_11520, n_11521, n_11522, a_SCH2ADDRREG_F2_G_aCLK, a_LC3_C2,
          a_EQ670, n_11526, n_11527, n_11528, n_11529, a_SCH0ADDRREG_F2_G,
          n_11531, n_11532, n_11533, n_11534, n_11535, n_11536, n_11537, n_11538,
          a_LC4_C2, a_EQ671, n_11541, n_11542, n_11543, n_11544, n_11545,
          n_11546, n_11547, n_11548, a_SCH0ADDRREG_F2_G_aCLRN, a_EQ869, n_11555,
          n_11556, n_11557, n_11558, n_11559, n_11560, n_11561, n_11562, n_11563,
          n_11564, n_11565, n_11566, n_11567, a_SCH0ADDRREG_F2_G_aCLK, a_N2543,
          a_EQ600, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576, n_11577,
          n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584, n_11585,
          n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592, n_11593,
          a_LC4_C11, a_EQ668, n_11596, n_11597, n_11598, n_11599, n_11600,
          n_11601, n_11602, a_SCH0ADDRREG_F3_G, n_11604, a_LC2_C11, a_EQ669,
          n_11607, n_11608, n_11609, n_11610, n_11611, n_11612, n_11613, n_11614,
          a_SCH0ADDRREG_F3_G_aCLRN, a_EQ870, n_11621, n_11622, n_11623, n_11624,
          n_11625, n_11626, n_11627, n_11628, n_11629, a_SCH0ADDRREG_F3_G_aCLK,
          a_LC3_C7, a_EQ286, n_11633, n_11634, n_11635, n_11636, n_11637,
          n_11638, n_11639, n_11640, n_11641, n_11642, n_11643, n_11644, n_11645,
          n_11646, n_11647, n_11648, n_11649, n_11650, n_11651, n_11652, n_11653,
          n_11654, a_LC4_C7, a_EQ719, n_11657, n_11658, n_11659, n_11660,
          n_11661, n_11662, n_11663, n_11664, n_11665, a_SCH2ADDRREG_F3_G,
          n_11667, a_SCH2ADDRREG_F3_G_aCLRN, a_EQ998, n_11674, n_11675, n_11676,
          n_11677, n_11678, n_11679, n_11680, n_11681, n_11682, n_11683, n_11684,
          n_11685, a_SCH2ADDRREG_F3_G_aCLK, a_LC4_C23, a_EQ693, n_11689, n_11690,
          n_11691, n_11692, n_11693, n_11694, n_11695, a_SCH1ADDRREG_F3_G,
          n_11697, a_LC5_C23, a_EQ694, n_11700, n_11701, n_11702, n_11703,
          n_11704, n_11705, n_11706, n_11707, a_SCH1ADDRREG_F3_G_aCLRN, a_EQ934,
          n_11714, n_11715, n_11716, n_11717, n_11718, n_11719, n_11720, n_11721,
          n_11722, a_SCH1ADDRREG_F3_G_aCLK, a_N944_aNOT, a_EQ329, n_11726,
          n_11727, n_11728, n_11729, n_11730, n_11731, n_11732, n_11733, n_11734,
          n_11735, n_11736, n_11737, n_11738, n_11739, n_11740, n_11741, n_11742,
          n_11743, n_11744, n_11745, n_11746, n_11747, a_LC3_C26, a_EQ745,
          n_11750, n_11751, n_11752, n_11753, n_11754, n_11755, n_11756, n_11757,
          n_11758, a_SCH3ADDRREG_F3_G, n_11760, a_SCH3ADDRREG_F3_G_aCLRN,
          a_EQ1062, n_11767, n_11768, n_11769, n_11770, n_11771, n_11772,
          n_11773, n_11774, n_11775, n_11776, a_SCH3ADDRREG_F3_G_aCLK, a_N2544,
          a_EQ601, n_11780, n_11781, n_11782, n_11783, n_11784, n_11785, n_11786,
          n_11787, n_11788, n_11789, n_11790, n_11791, n_11792, n_11793, n_11794,
          n_11795, n_11796, n_11797, n_11798, n_11799, n_11800, n_11801, n_11802,
          a_LC2_C23, a_EQ691, n_11805, n_11806, n_11807, n_11808, n_11809,
          n_11810, n_11811, a_SCH1ADDRREG_F4_G, n_11813, a_LC3_C23, a_EQ692,
          n_11816, n_11817, n_11818, n_11819, n_11820, n_11821, n_11822, n_11823,
          a_SCH1ADDRREG_F4_G_aCLRN, a_EQ935, n_11830, n_11831, n_11832, n_11833,
          n_11834, n_11835, n_11836, n_11837, n_11838, a_SCH1ADDRREG_F4_G_aCLK,
          a_LC6_C5, a_EQ287, n_11842, n_11843, n_11844, n_11845, n_11846,
          n_11847, n_11848, n_11849, n_11850, n_11851, n_11852, n_11853, n_11854,
          n_11855, n_11856, n_11857, n_11858, n_11859, n_11860, n_11861, n_11862,
          n_11863, a_LC3_C5, a_EQ718, n_11866, n_11867, n_11868, n_11869,
          n_11870, n_11871, n_11872, n_11873, n_11874, a_SCH2ADDRREG_F4_G,
          n_11876, a_SCH2ADDRREG_F4_G_aCLRN, a_EQ999, n_11883, n_11884, n_11885,
          n_11886, n_11887, n_11888, n_11889, n_11890, n_11891, n_11892, n_11893,
          n_11894, a_SCH2ADDRREG_F4_G_aCLK, a_N938_aNOT, a_EQ328, n_11898,
          n_11899, n_11900, n_11901, n_11902, n_11903, n_11904, n_11905, n_11906,
          n_11907, n_11908, n_11909, n_11910, n_11911, n_11912, n_11913, n_11914,
          n_11915, n_11916, n_11917, n_11918, n_11919, a_LC4_C1, a_EQ744,
          n_11922, n_11923, n_11924, n_11925, n_11926, n_11927, n_11928, n_11929,
          n_11930, a_SCH3ADDRREG_F4_G, n_11932, a_SCH3ADDRREG_F4_G_aCLRN,
          a_EQ1063, n_11939, n_11940, n_11941, n_11942, n_11943, n_11944,
          n_11945, n_11946, n_11947, n_11948, a_SCH3ADDRREG_F4_G_aCLK, a_LC6_C11,
          a_EQ666, n_11952, n_11953, n_11954, n_11955, n_11956, n_11957, n_11958,
          a_SCH0ADDRREG_F4_G, n_11960, a_LC5_C11, a_EQ667, n_11963, n_11964,
          n_11965, n_11966, n_11967, n_11968, n_11969, n_11970, a_SCH0ADDRREG_F4_G_aCLRN,
          a_EQ871, n_11977, n_11978, n_11979, n_11980, n_11981, n_11982, n_11983,
          n_11984, n_11985, a_SCH0ADDRREG_F4_G_aCLK, a_N2545, a_EQ602, n_11989,
          n_11990, n_11991, n_11992, n_11993, n_11994, n_11995, n_11996, n_11997,
          n_11998, n_11999, n_12000, n_12001, a_LC2_F23, a_EQ689, n_12004,
          n_12005, n_12006, n_12007, a_SCH1ADDRREG_F5_G, n_12009, n_12010,
          n_12011, n_12012, n_12013, n_12014, n_12015, n_12016, a_LC4_F23,
          a_EQ690, n_12019, n_12020, n_12021, n_12022, n_12023, n_12024, n_12025,
          n_12026, a_SCH1ADDRREG_F5_G_aCLRN, a_EQ936, n_12033, n_12034, n_12035,
          n_12036, n_12037, n_12038, n_12039, n_12040, n_12041, n_12042, n_12043,
          n_12044, n_12045, a_SCH1ADDRREG_F5_G_aCLK, a_LC3_F20, a_EQ716, n_12049,
          n_12050, n_12051, n_12052, n_12053, n_12054, n_12055, a_SCH2ADDRREG_F5_G,
          n_12057, a_LC1_F20, a_EQ717, n_12060, n_12061, n_12062, n_12063,
          n_12064, n_12065, n_12066, n_12067, n_12068, n_12069, n_12070, n_12071,
          n_12072, a_SCH2ADDRREG_F5_G_aCLRN, a_EQ1000, n_12079, n_12080, n_12081,
          n_12082, n_12083, n_12084, n_12085, n_12086, n_12087, a_SCH2ADDRREG_F5_G_aCLK,
          a_LC1_F21, a_EQ742, n_12091, n_12092, n_12093, n_12094, n_12095,
          n_12096, n_12097, n_12098, n_12099, a_SCH3ADDRREG_F5_G, n_12101,
          a_LC3_F21, a_EQ743, n_12104, n_12105, n_12106, n_12107, n_12108,
          n_12109, n_12110, a_SCH3ADDRREG_F5_G_aCLRN, a_EQ1064, n_12117, n_12118,
          n_12119, n_12120, n_12121, n_12122, n_12123, n_12124, n_12125, n_12126,
          n_12127, n_12128, n_12129, a_SCH3ADDRREG_F5_G_aCLK, a_LC3_F3, a_EQ664,
          n_12133, n_12134, n_12135, n_12136, a_SCH0ADDRREG_F5_G, n_12138,
          n_12139, n_12140, n_12141, n_12142, n_12143, n_12144, n_12145, a_LC4_F3,
          a_EQ665, n_12148, n_12149, n_12150, n_12151, n_12152, n_12153, n_12154,
          n_12155, a_SCH0ADDRREG_F5_G_aCLRN, a_EQ872, n_12162, n_12163, n_12164,
          n_12165, n_12166, n_12167, n_12168, n_12169, n_12170, n_12171, n_12172,
          n_12173, n_12174, a_SCH0ADDRREG_F5_G_aCLK, a_LC3_F14, a_EQ288, n_12178,
          n_12179, n_12180, n_12181, n_12182, n_12183, n_12184, n_12185, n_12186,
          n_12187, n_12188, n_12189, n_12190, n_12191, n_12192, n_12193, n_12194,
          n_12195, n_12196, n_12197, n_12198, n_12199, a_LC4_F14, a_EQ715,
          n_12202, n_12203, n_12204, n_12205, n_12206, n_12207, n_12208, n_12209,
          n_12210, a_SCH2ADDRREG_F6_G, n_12212, a_SCH2ADDRREG_F6_G_aCLRN,
          a_EQ1001, n_12219, n_12220, n_12221, n_12222, n_12223, n_12224,
          n_12225, n_12226, n_12227, n_12228, n_12229, n_12230, a_SCH2ADDRREG_F6_G_aCLK,
          a_N2546, a_EQ603, n_12234, n_12235, n_12236, n_12237, n_12238, n_12239,
          n_12240, n_12241, n_12242, n_12243, n_12244, n_12245, n_12246, n_12247,
          n_12248, n_12249, n_12250, n_12251, n_12252, n_12253, n_12254, n_12255,
          n_12256, a_LC5_F3, a_EQ662, n_12259, n_12260, n_12261, n_12262,
          a_SCH0ADDRREG_F6_G, n_12264, n_12265, n_12266, n_12267, n_12268,
          n_12269, n_12270, n_12271, a_LC2_F3, a_EQ663, n_12274, n_12275,
          n_12276, n_12277, n_12278, n_12279, n_12280, n_12281, a_SCH0ADDRREG_F6_G_aCLRN,
          a_EQ873, n_12288, n_12289, n_12290, n_12291, n_12292, n_12293, n_12294,
          n_12295, n_12296, n_12297, n_12298, n_12299, n_12300, a_SCH0ADDRREG_F6_G_aCLK,
          a_LC5_F23, a_EQ687, n_12304, n_12305, n_12306, n_12307, a_SCH1ADDRREG_F6_G,
          n_12309, n_12310, n_12311, n_12312, n_12313, n_12314, n_12315, n_12316,
          a_LC1_F23, a_EQ688, n_12319, n_12320, n_12321, n_12322, n_12323,
          n_12324, n_12325, n_12326, a_SCH1ADDRREG_F6_G_aCLRN, a_EQ937, n_12333,
          n_12334, n_12335, n_12336, n_12337, n_12338, n_12339, n_12340, n_12341,
          n_12342, n_12343, n_12344, n_12345, a_SCH1ADDRREG_F6_G_aCLK, a_N933_aNOT,
          a_EQ326, n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355,
          n_12356, n_12357, n_12358, n_12359, n_12360, n_12361, n_12362, n_12363,
          n_12364, n_12365, n_12366, n_12367, n_12368, n_12369, n_12370, a_LC4_F21,
          a_EQ741, n_12373, n_12374, n_12375, n_12376, n_12377, n_12378, n_12379,
          n_12380, n_12381, a_SCH3ADDRREG_F6_G, n_12383, a_SCH3ADDRREG_F6_G_aCLRN,
          a_EQ1065, n_12390, n_12391, n_12392, n_12393, n_12394, n_12395,
          n_12396, n_12397, n_12398, n_12399, a_SCH3ADDRREG_F6_G_aCLK, a_LC6_D25,
          a_EQ739, n_12403, n_12404, n_12405, n_12406, n_12407, n_12408, n_12409,
          n_12410, n_12411, a_SCH3ADDRREG_F7_G, n_12413, a_LC4_D25, a_EQ740,
          n_12416, n_12417, n_12418, n_12419, n_12420, n_12421, n_12422, a_SCH3ADDRREG_F7_G_aCLRN,
          a_EQ1066, n_12429, n_12430, n_12431, n_12432, n_12433, n_12434,
          n_12435, n_12436, n_12437, n_12438, n_12439, n_12440, n_12441, a_SCH3ADDRREG_F7_G_aCLK,
          a_N786_aNOT, a_EQ299, n_12445, n_12446, n_12447, n_12448, n_12449,
          n_12450, n_12451, a_SCH2ADDRREG_F7_G, n_12453, a_LC4_D17, a_EQ714,
          n_12456, n_12457, n_12458, n_12459, n_12460, n_12461, n_12462, n_12463,
          n_12464, n_12465, n_12466, n_12467, n_12468, a_SCH2ADDRREG_F7_G_aCLRN,
          a_EQ1002, n_12475, n_12476, n_12477, n_12478, n_12479, n_12480,
          n_12481, n_12482, n_12483, a_SCH2ADDRREG_F7_G_aCLK, a_N2547, a_EQ604,
          n_12487, n_12488, n_12489, n_12490, n_12491, n_12492, n_12493, n_12494,
          n_12495, n_12496, n_12497, n_12498, n_12499, n_12500, n_12501, n_12502,
          n_12503, n_12504, n_12505, n_12506, n_12507, n_12508, n_12509, a_N183_aNOT,
          a_EQ204, n_12512, n_12513, n_12514, n_12515, n_12516, n_12517, n_12518,
          n_12519, a_SCH0ADDRREG_F7_G, n_12521, n_12522, n_12523, n_12524,
          a_LC3_D9, a_EQ661, n_12527, n_12528, n_12529, n_12530, n_12531,
          n_12532, n_12533, n_12534, a_SCH0ADDRREG_F7_G_aCLRN, a_EQ874, n_12541,
          n_12542, n_12543, n_12544, n_12545, n_12546, n_12547, n_12548, n_12549,
          n_12550, n_12551, n_12552, n_12553, a_SCH0ADDRREG_F7_G_aCLK, a_LC5_D19,
          a_EQ685, n_12557, n_12558, n_12559, n_12560, n_12561, n_12562, n_12563,
          n_12564, a_SCH1ADDRREG_F7_G, n_12566, n_12567, n_12568, n_12569,
          a_LC3_D19, a_EQ686, n_12572, n_12573, n_12574, n_12575, n_12576,
          n_12577, n_12578, n_12579, a_SCH1ADDRREG_F7_G_aCLRN, a_EQ938, n_12586,
          n_12587, n_12588, n_12589, n_12590, n_12591, n_12592, n_12593, n_12594,
          n_12595, n_12596, n_12597, n_12598, a_SCH1ADDRREG_F7_G_aCLK, a_LC8_B25,
          a_EQ430, n_12602, n_12603, n_12604, n_12605, n_12606, n_12607, n_12608,
          n_12609, a_N1467, a_EQ448, n_12612, n_12613, n_12614, n_12615, n_12616,
          n_12617, n_12618, a_N820_aCLRN, a_EQ306, n_12625, n_12626, n_12627,
          n_12628, n_12629, n_12630, n_12631, n_12632, n_12633, n_12634, a_N820_aCLK,
          a_LC2_D4, a_EQ360, n_12638, n_12639, n_12640, n_12641, n_12642,
          n_12643, n_12644, n_12645, n_12646, n_12647, n_12648, n_12649, a_N1141,
          a_EQ367, n_12652, n_12653, n_12654, n_12655, n_12656, n_12657, n_12658,
          n_12659, a_LC1_D4, a_EQ366, n_12662, n_12663, n_12664, n_12665,
          n_12666, n_12667, n_12668, n_12669, a_LC4_D12, a_EQ369, n_12672,
          n_12673, n_12674, n_12675, n_12676, n_12677, n_12678, n_12679, a_LC3_D12,
          a_EQ368, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687, n_12688,
          n_12689, a_N3541_aCLRN, a_EQ837, n_12696, n_12697, n_12698, n_12699,
          n_12700, n_12701, n_12702, n_12703, n_12704, n_12705, n_12706, n_12707,
          a_N3541_aCLK, a_N2395, a_N2395_aIN, n_12711, n_12712, n_12713, n_12714,
          n_12715, n_12716, a_LC4_B13, a_EQ392, n_12719, n_12720, n_12721,
          n_12722, n_12723, n_12724, n_12725, n_12726, a_N4179, a_N4179_aD,
          n_12734, n_12735, n_12736, n_12737, n_12738, a_N4179_aCLK, a_N4183,
          a_N4183_aD, n_12746, n_12747, n_12748, n_12749, n_12750, a_N4183_aCLK,
          a_N59, a_EQ182, n_12754, n_12755, n_12756, n_12757, n_12758, n_12759,
          n_12760, n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, a_N4178,
          a_N4178_aD, n_12774, n_12775, n_12776, n_12777, n_12778, a_N4178_aCLK,
          a_N4182, a_N4182_aD, n_12786, n_12787, n_12788, n_12789, n_12790,
          a_N4182_aCLK, a_N2534, a_EQ594, n_12794, n_12795, n_12796, n_12797,
          n_12798, n_12799, n_12800, n_12801, n_12802, n_12803, n_12804, n_12805,
          a_LC3_B6, a_EQ596, n_12808, n_12809, n_12810, n_12811, n_12812,
          n_12813, n_12814, n_12815, a_LC4_E2, a_EQ474, n_12818, n_12819,
          n_12820, n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827,
          n_12828, n_12829, n_12830, n_12831, a_LC1_E2, a_EQ473, n_12834,
          n_12835, n_12836, n_12837, n_12838, n_12839, n_12840, n_12841, n_12842,
          n_12843, n_12844, n_12845, n_12846, n_12847, a_N4180, a_N4180_aD,
          n_12855, n_12856, n_12857, n_12858, n_12859, a_N4180_aCLK, a_N4184,
          a_N4184_aD, n_12867, n_12868, n_12869, n_12870, n_12871, a_N4184_aCLK,
          a_N2536, a_EQ595, n_12875, n_12876, n_12877, n_12878, n_12879, n_12880,
          n_12881, n_12882, n_12883, n_12884, n_12885, n_12886, a_N4181, a_N4181_aD,
          n_12894, n_12895, n_12896, n_12897, n_12898, a_N4181_aCLK, a_N4185,
          a_N4185_aD, n_12906, n_12907, n_12908, n_12909, n_12910, a_N4185_aCLK,
          a_N55, a_EQ180, n_12914, n_12915, n_12916, n_12917, n_12918, n_12919,
          n_12920, n_12921, n_12922, n_12923, n_12924, n_12925, n_12926, a_LC4_B16,
          a_EQ597, n_12929, n_12930, n_12931, n_12932, n_12933, n_12934, n_12935,
          n_12936, a_N1585_aNOT, a_EQ475, n_12939, n_12940, n_12941, n_12942,
          n_12943, n_12944, n_12945, n_12946, n_12947, n_12948, a_LC1_E15,
          a_EQ469, n_12951, n_12952, n_12953, n_12954, n_12955, n_12956, n_12957,
          n_12958, a_LC6_E26, a_EQ470, n_12961, n_12962, n_12963, n_12964,
          n_12965, n_12966, n_12967, n_12968, a_N1581_aNOT, a_EQ471, n_12971,
          n_12972, n_12973, n_12974, n_12975, n_12976, n_12977, n_12978, a_N2394,
          a_N2394_aIN, n_12981, n_12982, n_12983, n_12984, n_12985, n_12986,
          n_12987, a_N2369_aNOT, a_N2369_aNOT_aIN, n_12990, n_12991, n_12992,
          n_12993, n_12994, n_12995, n_12996, a_LC4_B3, a_EQ393, n_13000,
          n_13001, n_13002, n_13003, n_13004, n_13005, n_13006, n_13007, n_13008,
          n_13009, n_13010, a_N2359_aNOT, a_N2359_aNOT_aIN, n_13013, n_13014,
          n_13015, n_13016, n_13017, a_LC3_B16, a_EQ394, n_13020, n_13021,
          n_13022, n_13023, n_13024, n_13025, n_13026, n_13027, a_N1249, a_N1249_aIN,
          n_13030, n_13031, n_13032, n_13033, n_13034, n_13035, n_13036, a_LC3_B3,
          a_EQ395, n_13039, n_13040, n_13041, n_13042, n_13043, n_13044, n_13045,
          n_13046, n_13047, n_13048, a_N822_aCLRN, a_EQ308, n_13055, n_13056,
          n_13057, n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064,
          n_13065, n_13066, a_N822_aCLK, a_N1387, a_N1387_aIN, n_13070, n_13071,
          n_13072, n_13073, n_13074, n_13075, a_LC8_B13, a_EQ429, n_13078,
          n_13079, n_13080, n_13081, n_13082, n_13083, n_13084, n_13085, n_13086,
          a_N821_aCLRN, a_EQ307, n_13093, n_13094, n_13095, n_13096, n_13097,
          n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104, a_N821_aCLK,
          a_STEMPORARYREG_F4_G, a_STEMPORARYREG_F4_G_aCLRN, a_EQ1185, n_13113,
          n_13114, n_13115, n_13116, n_13117, n_13118, n_13119, n_13120, n_13121,
          n_13122, n_13123, a_STEMPORARYREG_F4_G_aCLK, a_SCOMMANDREG_F7_G,
          a_SCOMMANDREG_F7_G_aCLRN, a_EQ1130, n_13132, n_13133, n_13134, n_13135,
          n_13136, n_13137, n_13138, n_13139, n_13140, n_13141, n_13142, a_SCOMMANDREG_F7_G_aCLK,
          a_N2606, a_EQ648, n_13146, n_13147, n_13148, n_13149, n_13150, n_13151,
          a_LC2_B2, a_EQ543, n_13154, n_13155, n_13156, n_13157, n_13158,
          n_13159, n_13160, n_13161, n_13162, a_LC6_B2, a_EQ544, n_13165,
          n_13166, n_13167, n_13168, n_13169, n_13170, n_13171, n_13172, a_LC7_B2,
          a_EQ545, n_13175, n_13176, n_13177, n_13178, n_13179, n_13180, n_13181,
          n_13182, n_13183, a_LC5_B2, a_EQ542, n_13186, n_13187, n_13188,
          n_13189, n_13190, n_13191, n_13192, n_13193, a_LC4_B2, a_EQ546,
          n_13196, n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203,
          a_N4186, a_N4186_aD, n_13211, n_13212, n_13213, n_13214, n_13215,
          a_N4186_aCLK, a_N4187, a_N4187_aD, n_13223, n_13224, n_13225, n_13226,
          n_13227, a_N4187_aCLK, a_N4170_aNOT, a_EQ853, n_13231, n_13232,
          n_13233, n_13234, n_13235, n_13236, a_SCHANNEL_F1_G_aCLRN, a_EQ866,
          n_13243, n_13244, n_13245, n_13246, n_13247, n_13248, n_13249, n_13250,
          n_13251, n_13252, n_13253, a_SCHANNEL_F1_G_aCLK, a_LC8_B26, a_EQ547,
          n_13257, n_13258, n_13259, n_13260, n_13261, n_13262, n_13263, n_13264,
          n_13265, n_13266, a_LC7_B26_aNOT, a_LC7_B26_aNOT_aIN, n_13269, n_13270,
          n_13271, n_13272, n_13273, a_LC6_B26, a_EQ549, n_13276, n_13277,
          n_13278, n_13279, n_13280, n_13281, n_13282, n_13283, a_LC4_B26,
          a_EQ550, n_13286, n_13287, n_13288, n_13289, n_13290, n_13291, n_13292,
          n_13293, n_13294, n_13295, a_LC3_B26, a_EQ551, n_13298, n_13299,
          n_13300, n_13301, n_13302, n_13303, n_13304, n_13305, a_LC2_B26,
          a_EQ552, n_13308, n_13309, n_13310, n_13311, n_13312, n_13313, n_13314,
          n_13315, a_SCHANNEL_F0_G_aCLRN, a_EQ865, n_13322, n_13323, n_13324,
          n_13325, n_13326, n_13327, n_13328, n_13329, n_13330, n_13331, n_13332,
          a_SCHANNEL_F0_G_aCLK, startdma_aD, n_13339, n_13340, n_13341, n_13342,
          n_13343, startdma_aCLK, a_SCOMMANDREG_F5_G, a_SCOMMANDREG_F5_G_aCLRN,
          a_EQ1128, n_13352, n_13353, n_13354, n_13355, n_13356, n_13357,
          n_13358, n_13359, n_13360, n_13361, n_13362, a_SCOMMANDREG_F5_G_aCLK,
          a_LC6_B3, a_EQ529, n_13366, n_13367, n_13368, n_13369, n_13370,
          n_13371, n_13372, n_13373, n_13374, a_LC7_B16, a_LC7_B16_aIN, n_13377,
          n_13378, n_13379, n_13380, n_13381, n_13382, a_LC8_B16, a_EQ531,
          n_13385, n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392,
          n_13393, n_13394, a_LC1_B2, a_LC1_B2_aIN, n_13397, n_13398, n_13399,
          n_13400, n_13401, n_13402, a_N1381, a_EQ428, n_13405, n_13406, n_13407,
          n_13408, n_13409, n_13410, n_13411, n_13412, n_13413, n_13414, n_13415,
          a_LC7_B3, a_EQ532, n_13418, n_13419, n_13420, n_13421, n_13422,
          n_13423, n_13424, n_13425, n_13426, n_13427, a_LC2_F17, a_EQ526,
          n_13430, n_13431, n_13432, n_13433, n_13434, n_13435, n_13436, n_13437,
          n_13438, n_13439, a_LC1_F17, a_EQ527, n_13442, n_13443, n_13444,
          n_13445, n_13446, n_13447, n_13448, n_13449, n_13450, n_13451, a_LC6_F17,
          a_EQ524, n_13454, n_13455, n_13456, n_13457, n_13458, n_13459, n_13460,
          n_13461, n_13462, n_13463, a_LC4_F17, a_EQ525, n_13466, n_13467,
          n_13468, n_13469, n_13470, n_13471, n_13472, n_13473, n_13474, n_13475,
          a_LC5_F17, a_EQ528, n_13478, n_13479, n_13480, n_13481, n_13482,
          n_13483, n_13484, n_13485, n_13486, n_13487, n_13488, n_13489, n_13490,
          n_13491, a_N823_aCLRN, a_EQ309, n_13498, n_13499, n_13500, n_13501,
          n_13502, n_13503, n_13504, n_13505, n_13506, n_13507, a_N823_aCLK,
          a_LC1_D18, a_EQ450, n_13511, n_13512, n_13513, n_13514, n_13515,
          n_13516, n_13517, n_13518, a_LC4_D18, a_EQ453, n_13521, n_13522,
          n_13523, n_13524, n_13525, n_13526, n_13527, n_13528, n_13529, n_13530,
          n_13531, n_13532, n_13533, n_13534, n_13535, n_13536, n_13537, a_N1486,
          a_EQ454, n_13540, n_13541, n_13542, n_13543, n_13544, n_13545, n_13546,
          n_13547, a_N1471, a_EQ452, n_13550, n_13551, n_13552, n_13553, n_13554,
          n_13555, n_13556, n_13557, n_13558, n_13559, a_LC2_D18, a_EQ451,
          n_13562, n_13563, n_13564, n_13565, n_13566, n_13567, n_13568, n_13569,
          a_LC7_D18_aCLRN, a_EQ044, n_13576, n_13577, n_13578, n_13579, n_13580,
          n_13581, n_13582, n_13583, n_13584, n_13585, n_13586, n_13587, a_LC7_D18_aCLK,
          a_LC4_C17, a_EQ523, n_13591, n_13592, n_13593, n_13594, n_13595,
          n_13596, n_13597, n_13598, n_13599, n_13600, n_13601, n_13602, a_N1904,
          a_EQ519, n_13605, n_13606, n_13607, n_13608, n_13609, n_13610, n_13611,
          n_13612, a_LC5_C17, a_EQ522, n_13615, n_13616, n_13617, n_13618,
          n_13619, n_13620, n_13621, n_13622, a_LC2_C17, a_EQ521, n_13625,
          n_13626, n_13627, n_13628, n_13629, n_13630, n_13631, n_13632, a_LC1_C17,
          a_EQ520, n_13635, n_13636, n_13637, n_13638, n_13639, n_13640, n_13641,
          n_13642, a_LC7_C17_aCLRN, a_EQ043, n_13649, n_13650, n_13651, n_13652,
          n_13653, n_13654, n_13655, n_13656, n_13657, n_13658, n_13659, n_13660,
          a_LC7_C17_aCLK, a_N1337_aNOT, a_EQ424, n_13664, n_13665, n_13666,
          n_13667, n_13668, n_13669, n_13670, n_13671, a_N1321, a_EQ413, n_13674,
          n_13675, n_13676, n_13677, n_13678, n_13679, n_13680, n_13681, a_LC8_C16,
          a_EQ412, n_13684, n_13685, n_13686, n_13687, n_13688, n_13689, n_13690,
          n_13691, a_LC2_C16, a_EQ415, n_13694, n_13695, n_13696, n_13697,
          n_13698, n_13699, n_13700, n_13701, a_LC5_C16, a_EQ414, n_13704,
          n_13705, n_13706, n_13707, n_13708, n_13709, n_13710, n_13711, a_LC4_C16_aCLRN,
          a_EQ042, n_13718, n_13719, n_13720, n_13721, n_13722, n_13723, n_13724,
          n_13725, n_13726, n_13727, n_13728, n_13729, a_LC4_C16_aCLK, a_LC5_C24,
          a_EQ289, n_13733, n_13734, n_13735, n_13736, n_13737, n_13738, n_13739,
          n_13740, a_LC6_C24, a_EQ290, n_13743, n_13744, n_13745, n_13746,
          n_13747, n_13748, n_13749, n_13750, a_N725_aNOT, a_EQ291, n_13753,
          n_13754, n_13755, n_13756, n_13757, n_13758, n_13759, n_13760, a_LC4_C24,
          a_EQ293, n_13763, n_13764, n_13765, n_13766, n_13767, n_13768, n_13769,
          n_13770, a_LC3_C24, a_EQ292, n_13773, n_13774, n_13775, n_13776,
          n_13777, n_13778, n_13779, n_13780, a_LC2_C24_aCLRN, a_EQ041, n_13787,
          n_13788, n_13789, n_13790, n_13791, n_13792, n_13793, n_13794, n_13795,
          n_13796, n_13797, n_13798, a_LC2_C24_aCLK, a_N1725_aNOT, a_EQ495,
          n_13802, n_13803, n_13804, n_13805, n_13806, n_13807, n_13808, n_13809,
          a_N1729, a_EQ497, n_13812, n_13813, n_13814, n_13815, n_13816, n_13817,
          n_13818, n_13819, a_LC3_C15, a_EQ489, n_13822, n_13823, n_13824,
          n_13825, n_13826, n_13827, n_13828, n_13829, a_LC3_C16, a_EQ491,
          n_13832, n_13833, n_13834, n_13835, n_13836, n_13837, n_13838, n_13839,
          a_LC4_C22, a_EQ490, n_13842, n_13843, n_13844, n_13845, n_13846,
          n_13847, n_13848, n_13849, a_LC1_C16_aCLRN, a_EQ040, n_13856, n_13857,
          n_13858, n_13859, n_13860, n_13861, n_13862, n_13863, n_13864, n_13865,
          n_13866, n_13867, a_LC1_C16_aCLK, a_LC6_F6, a_EQ237, n_13871, n_13872,
          n_13873, n_13874, n_13875, n_13876, n_13877, n_13878, a_LC5_F6,
          a_EQ238, n_13881, n_13882, n_13883, n_13884, n_13885, n_13886, n_13887,
          n_13888, a_N423_aNOT, a_EQ241, n_13891, n_13892, n_13893, n_13894,
          n_13895, n_13896, n_13897, n_13898, n_13899, n_13900, n_13901, n_13902,
          a_LC2_F6, a_EQ240, n_13905, n_13906, n_13907, n_13908, n_13909,
          n_13910, n_13911, n_13912, a_LC1_F6, a_EQ239, n_13915, n_13916,
          n_13917, n_13918, n_13919, n_13920, n_13921, n_13922, a_LC3_F6_aCLRN,
          a_EQ039, n_13929, n_13930, n_13931, n_13932, n_13933, n_13934, n_13935,
          n_13936, n_13937, n_13938, n_13939, n_13940, a_LC3_F6_aCLK, a_N1726_aNOT,
          a_EQ496, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949, n_13950,
          n_13951, a_N1730, a_EQ498, n_13954, n_13955, n_13956, n_13957, n_13958,
          n_13959, n_13960, n_13961, a_LC6_F10, a_EQ492, n_13964, n_13965,
          n_13966, n_13967, n_13968, n_13969, n_13970, n_13971, n_13972, n_13973,
          n_13974, n_13975, a_LC2_F10, a_EQ494, n_13978, n_13979, n_13980,
          n_13981, n_13982, n_13983, n_13984, n_13985, a_LC3_F10, a_EQ493,
          n_13988, n_13989, n_13990, n_13991, n_13992, n_13993, n_13994, n_13995,
          a_LC4_F10_aCLRN, a_EQ038, n_14002, n_14003, n_14004, n_14005, n_14006,
          n_14007, n_14008, n_14009, n_14010, n_14011, n_14012, n_14013, a_LC4_F10_aCLK,
          a_LC4_D27, a_EQ200, n_14017, n_14018, n_14019, n_14020, n_14021,
          n_14022, n_14023, n_14024, a_LC3_D27, a_EQ201, n_14027, n_14028,
          n_14029, n_14030, n_14031, n_14032, n_14033, n_14034, a_N185_aNOT,
          a_EQ205, n_14037, n_14038, n_14039, n_14040, n_14041, n_14042, n_14043,
          n_14044, a_LC2_D27, a_EQ203, n_14047, n_14048, n_14049, n_14050,
          n_14051, n_14052, n_14053, n_14054, a_LC1_D27, a_EQ202, n_14057,
          n_14058, n_14059, n_14060, n_14061, n_14062, n_14063, n_14064, a_LC5_D27_aCLRN,
          a_EQ037, n_14071, n_14072, n_14073, n_14074, n_14075, n_14076, n_14077,
          n_14078, n_14079, n_14080, n_14081, n_14082, a_LC5_D27_aCLK, a_LC7_B10,
          a_EQ110, n_14086, n_14087, n_14088, n_14089, n_14090, n_14091, n_14092,
          n_14093, n_14094, n_14095, n_14096, a_EQ864, n_14098, n_14099, n_14100,
          n_14101, n_14102, n_14103, a_N2389, a_EQ571, n_14106, n_14107, n_14108,
          n_14109, n_14110, n_14111, a_LC3_B9, a_EQ121, n_14114, n_14115,
          n_14116, n_14117, n_14118, n_14119, n_14120, n_14121, a_LC5_D23,
          a_EQ111, n_14124, n_14125, n_14126, n_14127, n_14128, n_14129, n_14130,
          n_14131, a_LC2_F9, a_EQ112, n_14134, n_14135, n_14136, n_14137,
          n_14138, n_14139, n_14140, n_14141, a_LC4_D23, a_EQ113, n_14144,
          n_14145, n_14146, n_14147, n_14148, n_14149, n_14150, n_14151, a_LC3_D23,
          a_EQ114, n_14154, n_14155, n_14156, n_14157, n_14158, n_14159, a_N2351,
          n_14161, n_14162, a_LC1_D23, a_EQ115, n_14165, n_14166, n_14167,
          n_14168, n_14169, n_14170, n_14171, n_14172, n_14173, n_14174, a_LC6_D22,
          a_EQ116, n_14177, n_14178, n_14179, n_14180, n_14181, n_14182, n_14183,
          n_14184, a_LC4_D22, a_EQ117, n_14187, n_14188, n_14189, n_14190,
          n_14191, n_14192, n_14193, n_14194, a_LC2_D22, a_EQ118, n_14197,
          n_14198, n_14199, n_14200, n_14201, n_14202, n_14203, n_14204, a_LC1_D22,
          a_EQ119, n_14207, n_14208, n_14209, n_14210, n_14211, n_14212, n_14213,
          n_14214, a_LC5_D22, a_EQ120, n_14217, n_14218, n_14219, n_14220,
          n_14221, n_14222, n_14223, n_14224, n_14225, n_14226, a_LC2_D23,
          a_EQ122, n_14229, n_14230, n_14231, n_14232, n_14233, n_14234, n_14235,
          n_14236, n_14237, n_14238, a_N1830, a_N1830_aIN, n_14241, n_14242,
          n_14243, n_14244, a_LC6_B10, a_EQ123, n_14247, n_14248, n_14249,
          n_14250, n_14251, n_14252, n_14253, n_14254, a_LC4_B10, a_EQ124,
          n_14257, n_14258, n_14259, n_14260, n_14261, n_14262, n_14263, n_14264,
          n_14265, a_EQ125, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272,
          n_14273, n_14274, n_14275, n_14276, n_14277, a_LC2_B21, a_EQ143,
          n_14280, n_14281, n_14282, n_14283, n_14284, n_14285, n_14286, n_14287,
          n_14288, n_14289, n_14290, a_LC8_C8, a_EQ152, n_14293, n_14294,
          n_14295, n_14296, n_14297, n_14298, n_14299, n_14300, a_LC7_C8,
          a_EQ153, n_14303, n_14304, n_14305, n_14306, n_14307, n_14308, n_14309,
          n_14310, a_LC5_C8, a_EQ154, n_14313, n_14314, n_14315, n_14316,
          n_14317, n_14318, n_14319, n_14320, a_LC4_C8, a_EQ155, n_14323,
          n_14324, n_14325, n_14326, n_14327, n_14328, n_14329, n_14330, a_LC6_C8,
          a_EQ156, n_14333, n_14334, n_14335, n_14336, n_14337, n_14338, n_14339,
          n_14340, n_14341, n_14342, a_LC4_A17, a_EQ148, n_14345, n_14346,
          n_14347, n_14348, n_14349, n_14350, n_14351, n_14352, a_LC3_A17,
          a_EQ149, n_14355, n_14356, n_14357, n_14358, n_14359, n_14360, n_14361,
          n_14362, a_LC2_A17, a_EQ150, n_14365, n_14366, n_14367, n_14368,
          n_14369, n_14370, n_14371, n_14372, a_LC1_A17, a_EQ151, n_14375,
          n_14376, n_14377, n_14378, n_14379, n_14380, n_14381, n_14382, a_LC5_A17,
          a_EQ147, n_14385, n_14386, n_14387, n_14388, n_14389, n_14390, n_14391,
          n_14392, a_LC6_A17, a_EQ157, n_14395, n_14396, n_14397, n_14398,
          n_14399, n_14400, n_14401, n_14402, n_14403, n_14404, n_14405, a_LC5_B23,
          a_EQ145, n_14408, n_14409, n_14410, n_14411, n_14412, n_14413, n_14414,
          n_14415, a_LC5_B21, a_EQ146, n_14418, n_14419, n_14420, n_14421,
          n_14422, n_14423, n_14424, n_14425, n_14426, a_LC4_B21, a_EQ144,
          n_14429, n_14430, n_14431, n_14432, n_14433, n_14434, n_14435, n_14436,
          a_LC7_B21, a_EQ158, n_14439, n_14440, n_14441, n_14442, n_14443,
          n_14444, n_14445, n_14446, a_EQ159, n_14448, n_14449, n_14450, n_14451,
          n_14452, n_14453, n_14454, n_14455, n_14456, n_14457, n_14458, n_14459,
          a_LC7_E23, a_EQ077, n_14462, n_14463, n_14464, n_14465, n_14466,
          n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, a_LC8_E26,
          a_EQ480, n_14475, n_14476, n_14477, n_14478, n_14479, n_14480, n_14481,
          n_14482, n_14483, n_14484, a_LC7_E26, a_EQ481, n_14487, n_14488,
          n_14489, n_14490, n_14491, n_14492, n_14493, n_14494, n_14495, n_14496,
          a_N1647_aNOT, a_EQ482, n_14499, n_14500, n_14501, n_14502, n_14503,
          n_14504, n_14505, n_14506, a_LC6_B7, a_EQ090, n_14509, n_14510,
          n_14511, n_14512, n_14513, n_14514, n_14515, n_14516, a_LC8_E23,
          a_EQ091, n_14519, n_14520, n_14521, n_14522, n_14523, n_14524, n_14525,
          n_14526, n_14527, a_LC4_B14, a_EQ088, n_14530, n_14531, n_14532,
          n_14533, n_14534, n_14535, n_14536, n_14537, a_LC2_C21, a_EQ078,
          n_14540, n_14541, n_14542, n_14543, n_14544, n_14545, n_14546, n_14547,
          a_LC7_C21, a_EQ079, n_14550, n_14551, n_14552, n_14553, n_14554,
          n_14555, n_14556, n_14557, a_LC6_C21, a_EQ080, n_14560, n_14561,
          n_14562, n_14563, n_14564, n_14565, n_14566, n_14567, a_LC4_C21,
          a_EQ081, n_14570, n_14571, n_14572, n_14573, n_14574, n_14575, n_14576,
          n_14577, a_LC5_C21, a_EQ082, n_14580, n_14581, n_14582, n_14583,
          n_14584, n_14585, n_14586, n_14587, n_14588, n_14589, a_LC5_E4,
          a_EQ083, n_14592, n_14593, n_14594, n_14595, n_14596, n_14597, n_14598,
          n_14599, a_LC4_E4, a_EQ084, n_14602, n_14603, n_14604, n_14605,
          n_14606, n_14607, n_14608, n_14609, a_LC4_E27, a_EQ085, n_14612,
          n_14613, n_14614, n_14615, n_14616, n_14617, n_14618, n_14619, a_LC2_E18,
          a_EQ086, n_14622, n_14623, n_14624, n_14625, n_14626, n_14627, n_14628,
          n_14629, a_LC3_E4, a_EQ087, n_14632, n_14633, n_14634, n_14635,
          n_14636, n_14637, n_14638, n_14639, n_14640, n_14641, a_LC6_E4,
          a_EQ089, n_14644, n_14645, n_14646, n_14647, n_14648, n_14649, n_14650,
          n_14651, n_14652, n_14653, a_EQ092, n_14655, n_14656, n_14657, n_14658,
          n_14659, n_14660, n_14661, n_14662, n_14663, n_14664, n_14665, a_LC2_A27,
          a_EQ060, n_14668, n_14669, n_14670, n_14671, n_14672, n_14673, n_14674,
          n_14675, a_LC6_A10, a_EQ066, n_14678, n_14679, n_14680, n_14681,
          n_14682, n_14683, n_14684, n_14685, a_LC5_A10, a_EQ067, n_14688,
          n_14689, n_14690, n_14691, n_14692, n_14693, n_14694, n_14695, a_LC4_A10,
          a_EQ068, n_14698, n_14699, n_14700, n_14701, n_14702, n_14703, n_14704,
          n_14705, a_LC3_A10, a_EQ069, n_14708, n_14709, n_14710, n_14711,
          n_14712, n_14713, n_14714, n_14715, a_LC1_A10, a_EQ070, n_14718,
          n_14719, n_14720, n_14721, n_14722, n_14723, n_14724, n_14725, n_14726,
          n_14727, a_LC6_C13, a_EQ062, n_14730, n_14731, n_14732, n_14733,
          n_14734, n_14735, n_14736, n_14737, a_LC3_C8, a_EQ063, n_14740,
          n_14741, n_14742, n_14743, n_14744, n_14745, n_14746, n_14747, a_LC2_C8,
          a_EQ064, n_14750, n_14751, n_14752, n_14753, n_14754, n_14755, n_14756,
          n_14757, a_LC1_C8, a_EQ065, n_14760, n_14761, n_14762, n_14763,
          n_14764, n_14765, n_14766, n_14767, a_LC8_C19, a_EQ061, n_14770,
          n_14771, n_14772, n_14773, n_14774, n_14775, n_14776, n_14777, a_LC2_A10,
          a_EQ071, n_14780, n_14781, n_14782, n_14783, n_14784, n_14785, n_14786,
          n_14787, n_14788, n_14789, n_14790, a_LC1_A27, a_EQ072, n_14793,
          n_14794, n_14795, n_14796, n_14797, n_14798, n_14799, a_LC5_E10,
          a_EQ484, n_14802, n_14803, n_14804, n_14805, n_14806, n_14807, n_14808,
          n_14809, n_14810, n_14811, a_LC7_E10, a_EQ485, n_14814, n_14815,
          n_14816, n_14817, n_14818, n_14819, n_14820, n_14821, n_14822, n_14823,
          a_N1671_aNOT, a_EQ483, n_14826, n_14827, n_14828, n_14829, n_14830,
          n_14831, n_14832, n_14833, a_LC4_B7, a_EQ073, n_14836, n_14837,
          n_14838, n_14839, n_14840, n_14841, n_14842, n_14843, a_LC2_B18,
          a_EQ074, n_14846, n_14847, n_14848, n_14849, n_14850, n_14851, n_14852,
          n_14853, a_LC6_B18, a_EQ075, n_14856, n_14857, n_14858, n_14859,
          n_14860, n_14861, n_14862, n_14863, a_EQ076, n_14865, n_14866, n_14867,
          n_14868, n_14869, n_14870, n_14871, n_14872, n_14873, n_14874, n_14875,
          a_LC8_A27, a_EQ139, n_14878, n_14879, n_14880, n_14881, n_14882,
          n_14883, n_14884, n_14885, n_14886, n_14887, a_LC5_B7, a_EQ389,
          n_14890, n_14891, n_14892, n_14893, n_14894, n_14895, n_14896, n_14897,
          a_LC6_B27, a_EQ486, n_14900, n_14901, n_14902, n_14903, n_14904,
          n_14905, n_14906, n_14907, n_14908, n_14909, a_LC5_B27, a_EQ487,
          n_14912, n_14913, n_14914, n_14915, n_14916, n_14917, n_14918, n_14919,
          n_14920, n_14921, a_N1693_aNOT, a_EQ488, n_14924, n_14925, n_14926,
          n_14927, n_14928, n_14929, n_14930, n_14931, a_LC1_B27, a_EQ140,
          n_14934, n_14935, n_14936, n_14937, n_14938, n_14939, n_14940, a_LC8_B14,
          a_EQ137, n_14943, n_14944, n_14945, n_14946, n_14947, n_14948, n_14949,
          n_14950, n_14951, n_14952, a_LC1_C19, a_EQ127, n_14955, n_14956,
          n_14957, n_14958, n_14959, n_14960, n_14961, n_14962, a_LC4_C19,
          a_EQ128, n_14965, n_14966, n_14967, n_14968, n_14969, n_14970, n_14971,
          n_14972, a_LC5_C19, a_EQ129, n_14975, n_14976, n_14977, n_14978,
          n_14979, n_14980, n_14981, n_14982, a_LC6_C19, a_EQ130, n_14985,
          n_14986, n_14987, n_14988, n_14989, n_14990, n_14991, n_14992, a_LC2_C19,
          a_EQ131, n_14995, n_14996, n_14997, n_14998, n_14999, n_15000, n_15001,
          n_15002, n_15003, n_15004, a_LC6_A6, a_EQ132, n_15007, n_15008,
          n_15009, n_15010, n_15011, n_15012, n_15013, n_15014, a_LC5_A6,
          a_EQ133, n_15017, n_15018, n_15019, n_15020, n_15021, n_15022, n_15023,
          n_15024, a_LC4_A6, a_EQ134, n_15027, n_15028, n_15029, n_15030,
          n_15031, n_15032, n_15033, n_15034, a_LC3_A6, a_EQ135, n_15037,
          n_15038, n_15039, n_15040, n_15041, n_15042, n_15043, n_15044, a_LC2_A6,
          a_EQ136, n_15047, n_15048, n_15049, n_15050, n_15051, n_15052, n_15053,
          n_15054, n_15055, n_15056, a_LC1_A6, a_EQ138, n_15059, n_15060,
          n_15061, n_15062, n_15063, n_15064, n_15065, n_15066, n_15067, n_15068,
          a_LC7_A27, a_EQ141, n_15071, n_15072, n_15073, n_15074, n_15075,
          n_15076, n_15077, n_15078, n_15079, n_15080, n_15081, a_LC6_A27,
          a_EQ126, n_15084, n_15085, n_15086, n_15087, n_15088, n_15089, n_15090,
          n_15091, a_EQ142, n_15093, n_15094, n_15095, n_15096, n_15097, n_15098,
          n_15099, n_15100, a_LC6_E1, a_EQ510, n_15103, n_15104, n_15105,
          n_15106, n_15107, n_15108, n_15109, n_15110, n_15111, n_15112, a_LC5_E1,
          a_EQ511, n_15115, n_15116, n_15117, n_15118, n_15119, n_15120, n_15121,
          n_15122, n_15123, n_15124, a_N1837_aNOT, a_EQ509, n_15127, n_15128,
          n_15129, n_15130, n_15131, n_15132, n_15133, n_15134, a_LC8_F11,
          a_EQ095, n_15137, n_15138, n_15139, n_15140, n_15141, n_15142, n_15143,
          n_15144, a_LC7_F11, a_EQ096, n_15147, n_15148, n_15149, n_15150,
          n_15151, n_15152, n_15153, n_15154, a_LC6_F19, a_EQ097, n_15157,
          n_15158, n_15159, n_15160, n_15161, n_15162, n_15163, n_15164, a_LC6_F11,
          a_EQ098, n_15167, n_15168, n_15169, n_15170, n_15171, n_15172, n_15173,
          n_15174, a_LC3_F11, a_EQ099, n_15177, n_15178, n_15179, n_15180,
          n_15181, n_15182, n_15183, n_15184, n_15185, n_15186, a_LC7_E7,
          a_EQ100, n_15189, n_15190, n_15191, n_15192, n_15193, n_15194, n_15195,
          n_15196, a_LC6_E7, a_EQ101, n_15199, n_15200, n_15201, n_15202,
          n_15203, n_15204, n_15205, n_15206, a_LC5_E7, a_EQ102, n_15209,
          n_15210, n_15211, n_15212, n_15213, n_15214, n_15215, n_15216, a_LC2_E14,
          a_EQ103, n_15219, n_15220, n_15221, n_15222, n_15223, n_15224, n_15225,
          n_15226, a_LC4_E7, a_EQ104, n_15229, n_15230, n_15231, n_15232,
          n_15233, n_15234, n_15235, n_15236, n_15237, n_15238, a_LC3_E7,
          a_EQ105, n_15241, n_15242, n_15243, n_15244, n_15245, n_15246, n_15247,
          n_15248, n_15249, n_15250, a_N1849, a_N1849_aIN, n_15253, n_15254,
          n_15255, n_15256, n_15257, a_LC2_E7, a_EQ106, n_15260, n_15261,
          n_15262, n_15263, n_15264, n_15265, n_15266, n_15267, n_15268, a_LC6_B24,
          a_EQ107, n_15271, n_15272, n_15273, n_15274, n_15275, n_15276, n_15277,
          n_15278, a_LC2_B24, a_EQ108, n_15281, n_15282, n_15283, n_15284,
          n_15285, n_15286, n_15287, n_15288, n_15289, n_15290, n_15291, n_15292,
          a_EQ109, n_15294, n_15295, n_15296, n_15297, n_15298, n_15299, n_15300,
          n_15301, n_15302, n_15303, n_15304, a_LC5_B14, a_EQ055, n_15307,
          n_15308, n_15309, n_15310, n_15311, n_15312, n_15313, n_15314, n_15315,
          n_15316, n_15317, n_15318, n_15319, a_LC7_E18, a_EQ045, n_15322,
          n_15323, n_15324, n_15325, n_15326, n_15327, n_15328, n_15329, a_LC7_F19,
          a_EQ046, n_15332, n_15333, n_15334, n_15335, n_15336, n_15337, n_15338,
          n_15339, a_LC6_E18, a_EQ047, n_15342, n_15343, n_15344, n_15345,
          n_15346, n_15347, n_15348, n_15349, a_LC5_E18, a_EQ048, n_15352,
          n_15353, n_15354, n_15355, n_15356, n_15357, n_15358, n_15359, a_LC4_E18,
          a_EQ049, n_15362, n_15363, n_15364, n_15365, n_15366, n_15367, n_15368,
          n_15369, n_15370, n_15371, a_LC5_F11, a_EQ050, n_15374, n_15375,
          n_15376, n_15377, n_15378, n_15379, n_15380, n_15381, a_LC3_F26,
          a_EQ051, n_15384, n_15385, n_15386, n_15387, n_15388, n_15389, n_15390,
          n_15391, a_LC4_F11, a_EQ052, n_15394, n_15395, n_15396, n_15397,
          n_15398, n_15399, n_15400, n_15401, a_LC2_F11, a_EQ053, n_15404,
          n_15405, n_15406, n_15407, n_15408, n_15409, n_15410, n_15411, a_LC1_F11,
          a_EQ054, n_15414, n_15415, n_15416, n_15417, n_15418, n_15419, n_15420,
          n_15421, n_15422, n_15423, a_LC3_E18, a_EQ056, n_15426, n_15427,
          n_15428, n_15429, n_15430, n_15431, n_15432, n_15433, n_15434, n_15435,
          a_LC8_E2, a_EQ499, n_15438, n_15439, n_15440, n_15441, n_15442,
          n_15443, n_15444, n_15445, n_15446, n_15447, a_LC7_E2, a_EQ500,
          n_15450, n_15451, n_15452, n_15453, n_15454, n_15455, n_15456, n_15457,
          n_15458, n_15459, a_N1742_aNOT, a_EQ501, n_15462, n_15463, n_15464,
          n_15465, n_15466, n_15467, n_15468, n_15469, a_LC4_E23, a_EQ057,
          n_15472, n_15473, n_15474, n_15475, n_15476, n_15477, n_15478, n_15479,
          n_15480, a_LC3_E23, a_EQ058, n_15483, n_15484, n_15485, n_15486,
          n_15487, n_15488, n_15489, n_15490, n_15491, n_15492, n_15493, a_EQ059,
          n_15495, n_15496, n_15497, n_15498, n_15499, n_15500, n_15501, n_15502,
          n_15503, n_15504, n_15505, n_15506, n_15507, n_15508, a_N565_aNOT,
          a_EQ269, n_15511, n_15512, n_15513, n_15514, n_15515, n_15516, n_15517,
          n_15518, n_15519, n_15520, a_LC8_D15, a_EQ161, n_15523, n_15524,
          n_15525, n_15526, n_15527, n_15528, n_15529, n_15530, a_LC7_D15,
          a_EQ162, n_15533, n_15534, n_15535, n_15536, n_15537, n_15538, n_15539,
          n_15540, a_LC6_D15, a_EQ163, n_15543, n_15544, n_15545, n_15546,
          n_15547, n_15548, n_15549, n_15550, a_LC5_D15, a_EQ164, n_15553,
          n_15554, n_15555, n_15556, n_15557, n_15558, n_15559, n_15560, a_LC3_D15,
          a_EQ165, n_15563, n_15564, n_15565, n_15566, n_15567, n_15568, n_15569,
          n_15570, n_15571, n_15572, a_LC6_D13, a_EQ166, n_15575, n_15576,
          n_15577, n_15578, n_15579, n_15580, n_15581, n_15582, a_LC5_D13,
          a_EQ167, n_15585, n_15586, n_15587, n_15588, n_15589, n_15590, n_15591,
          n_15592, a_LC4_D13, a_EQ168, n_15595, n_15596, n_15597, n_15598,
          n_15599, n_15600, n_15601, n_15602, a_LC2_D13, a_EQ169, n_15605,
          n_15606, n_15607, n_15608, n_15609, n_15610, n_15611, n_15612, a_LC1_D13,
          a_EQ170, n_15615, n_15616, n_15617, n_15618, n_15619, n_15620, n_15621,
          n_15622, n_15623, n_15624, a_LC3_D13, a_EQ171, n_15627, n_15628,
          n_15629, n_15630, n_15631, n_15632, n_15633, n_15634, n_15635, n_15636,
          a_N1226_aNOT, a_N1226_aNOT_aIN, n_15639, n_15640, n_15641, n_15642,
          n_15643, a_LC6_E24, a_EQ160, n_15646, n_15647, n_15648, n_15649,
          n_15650, n_15651, n_15652, n_15653, n_15654, a_LC2_E24, a_EQ172,
          n_15657, n_15658, n_15659, n_15660, n_15661, n_15662, n_15663, n_15664,
          a_LC7_E15, a_EQ387, n_15667, n_15668, n_15669, n_15670, n_15671,
          n_15672, n_15673, n_15674, n_15675, n_15676, a_LC3_E26, a_EQ388,
          n_15679, n_15680, n_15681, n_15682, n_15683, n_15684, n_15685, n_15686,
          n_15687, n_15688, a_LC1_E24, a_EQ173, n_15691, n_15692, n_15693,
          n_15694, n_15695, n_15696, n_15697, n_15698, n_15699, n_15700, a_EQ174,
          n_15702, n_15703, n_15704, n_15705, n_15706, n_15707, n_15708, n_15709,
          n_15710, n_15711, n_15712, a_N2588, a_EQ641, n_15715, n_15716, n_15717,
          n_15718, n_15719, n_15720, n_15721, n_15722, n_15723, n_15724, n_15725,
          a_EQ094, n_15727, n_15728, n_15729, n_15730, n_15731, n_15732, n_15733,
          n_15734, n_15735, n_15736, n_15737, n_15738, n_15739, n_15740, n_15741,
          n_15742, a_EQ093, n_15744, n_15745, n_15746, n_15747, n_15748, n_15749,
          n_15750, n_15751, n_15752, n_15753, n_15754, n_15755, n_15756, n_15757,
          n_15758, n_15759, a_EQ176, n_15761, n_15762, n_15763, n_15764, n_15765,
          n_15766, n_15767, n_15768, n_15769, n_15770, n_15771, n_15772, n_15773,
          n_15774, n_15775, n_15776, a_EQ175, n_15778, n_15779, n_15780, n_15781,
          n_15782, n_15783, n_15784, n_15785, n_15786, n_15787, n_15788, n_15789,
          n_15790, n_15791, n_15792, n_15793, a_N2400, a_EQ578, n_15796, n_15797,
          n_15798, n_15799, n_15800, n_15801, n_15802, n_15803, n_15804, n_15805,
          a_LC5_B5, a_EQ1172, n_15808, n_15809, n_15810, n_15811, n_15812,
          n_15813, n_15814, n_15815, a_N2368, a_EQ564, n_15818, n_15819, n_15820,
          n_15821, n_15822, n_15823, n_15824, n_15825, n_15826, a_LC7_B5,
          a_EQ1171, n_15829, n_15830, n_15831, n_15832, n_15833, n_15834,
          n_15835, n_15836, n_15837, a_LC2_B5, a_EQ447, n_15840, n_15841,
          n_15842, n_15843, n_15844, n_15845, n_15846, n_15847, n_15848, n_15849,
          n_15850, a_N1468, a_EQ449, n_15853, n_15854, n_15855, n_15856, n_15857,
          n_15858, n_15859, n_15860, n_15861, n_15862, a_EQ1170, n_15864,
          n_15865, n_15866, n_15867, n_15868, n_15869, n_15870, n_15871, n_15872,
          a_LC5_B25, a_EQ1168, n_15875, n_15876, n_15877, n_15878, n_15879,
          n_15880, n_15881, n_15882, n_15883, n_15884, a_EQ1167, n_15886,
          n_15887, n_15888, n_15889, n_15890, n_15891, n_15892, n_15893, n_15894,
          a_LC2_B20, a_EQ1166, n_15897, n_15898, n_15899, n_15900, n_15901,
          n_15902, n_15903, n_15904, n_15905, n_15906, a_EQ1165, n_15908,
          n_15909, n_15910, n_15911, n_15912, n_15913, n_15914, n_15915, n_15916,
          a_N1252, a_EQ396, n_15919, n_15920, n_15921, n_15922, n_15923, n_15924,
          n_15925, n_15926, n_15927, n_15928, n_15929, n_15930, n_15931, n_15932,
          n_15933, n_15934, a_EQ1131, n_15936, n_15937, n_15938, n_15939,
          n_15940, n_15941, n_15942, n_15943, a_LC6_B16_aNOT_aIN, n_15945,
          n_15946, n_15947, n_15948, n_15949, n_15950, a_N2370_aNOT, a_N2370_aNOT_aIN,
          n_15953, n_15954, n_15955, n_15956, n_15957, n_15958, a_EQ862, n_15960,
          n_15961, n_15962, n_15963, n_15964, n_15965, n_15966, n_15967, n_15968,
          n_15969, n_15970, a_EQ196, n_15972, n_15973, n_15974, n_15975, n_15976,
          n_15977, a_EQ633, n_15979, n_15980, n_15981, n_15982, n_15983, n_15984,
          a_EQ555, n_15986, n_15987, n_15988, n_15989, n_15990, n_15991, n_15992,
          n_15993, n_15994, n_15995, a_EQ628, n_15997, n_15998, n_15999, n_16000,
          n_16001, n_16002, a_SCH1BWORDOUT_F1_G_aCLRN, a_EQ964, n_16009, n_16010,
          n_16011, n_16012, n_16013, n_16014, n_16015, n_16016, n_16017, a_SCH1BWORDOUT_F1_G_aCLK,
          a_EQ635, n_16020, n_16021, n_16022, n_16023, n_16024, n_16025, a_EQ629,
          n_16027, n_16028, n_16029, n_16030, n_16031, n_16032, a_SCH1BWORDOUT_F9_G_aCLRN,
          a_EQ972, n_16039, n_16040, n_16041, n_16042, n_16043, n_16044, n_16045,
          n_16046, n_16047, a_SCH1BWORDOUT_F9_G_aCLK, a_SCH1BWORDOUT_F10_G_aCLRN,
          a_EQ973, n_16055, n_16056, n_16057, n_16058, n_16059, n_16060, n_16061,
          n_16062, n_16063, a_SCH1BWORDOUT_F10_G_aCLK, a_EQ553, n_16066, n_16067,
          n_16068, n_16069, n_16070, n_16071, n_16072, n_16073, n_16074, n_16075,
          a_EQ625, n_16077, n_16078, n_16079, n_16080, n_16081, n_16082, n_16083,
          n_16084, a_SCH3BWORDOUT_F6_G_aCLRN, a_EQ1097, n_16091, n_16092,
          n_16093, n_16094, n_16095, n_16096, n_16097, n_16098, n_16099, a_SCH3BWORDOUT_F6_G_aCLK,
          a_SCH3BWORDOUT_F1_G_aCLRN, a_EQ1092, n_16107, n_16108, n_16109,
          n_16110, n_16111, n_16112, n_16113, n_16114, n_16115, a_SCH3BWORDOUT_F1_G_aCLK,
          a_EQ183, n_16118, n_16119, n_16120, n_16121, n_16122, n_16123, n_16124,
          n_16125, n_16126, n_16127, a_EQ627, n_16129, n_16130, n_16131, n_16132,
          n_16133, n_16134, a_SCH2BWORDOUT_F1_G_aCLRN, a_EQ1028, n_16141,
          n_16142, n_16143, n_16144, n_16145, n_16146, n_16147, n_16148, n_16149,
          a_SCH2BWORDOUT_F1_G_aCLK, a_SCH1BWORDOUT_F0_G_aCLRN, a_EQ963, n_16157,
          n_16158, n_16159, n_16160, n_16161, n_16162, n_16163, n_16164, n_16165,
          a_SCH1BWORDOUT_F0_G_aCLK, a_EQ557, n_16168, n_16169, n_16170, n_16171,
          n_16172, n_16173, n_16174, n_16175, n_16176, n_16177, a_EQ630, n_16179,
          n_16180, n_16181, n_16182, n_16183, n_16184, a_SCH0BWORDOUT_F1_G_aCLRN,
          a_EQ900, n_16191, n_16192, n_16193, n_16194, n_16195, n_16196, n_16197,
          n_16198, n_16199, a_SCH0BWORDOUT_F1_G_aCLK, a_SCH0BWORDOUT_F9_G_aCLRN,
          a_EQ908, n_16207, n_16208, n_16209, n_16210, n_16211, n_16212, n_16213,
          n_16214, n_16215, n_16216, n_16217, n_16218, n_16219, a_SCH0BWORDOUT_F9_G_aCLK,
          a_SCH2BWORDOUT_F9_G_aCLRN, a_EQ1036, n_16227, n_16228, n_16229,
          n_16230, n_16231, n_16232, n_16233, n_16234, n_16235, n_16236, n_16237,
          n_16238, n_16239, a_SCH2BWORDOUT_F9_G_aCLK, a_SCH1BWORDOUT_F2_G_aCLRN,
          a_EQ965, n_16247, n_16248, n_16249, n_16250, n_16251, n_16252, n_16253,
          n_16254, n_16255, a_SCH1BWORDOUT_F2_G_aCLK, a_SCH0BWORDOUT_F3_G_aCLRN,
          a_EQ902, n_16263, n_16264, n_16265, n_16266, n_16267, n_16268, n_16269,
          n_16270, n_16271, a_SCH0BWORDOUT_F3_G_aCLK, a_SCH1BWORDOUT_F3_G_aCLRN,
          a_EQ966, n_16279, n_16280, n_16281, n_16282, n_16283, n_16284, n_16285,
          n_16286, n_16287, a_SCH1BWORDOUT_F3_G_aCLK : std_logic;

COMPONENT TRIBUF_a8237
    PORT (in1, oe  : IN std_logic; y : OUT std_logic);
END COMPONENT;

COMPONENT DFF_a8237
    PORT (d, clk, clrn, prn : IN std_logic; q : OUT std_logic);
END COMPONENT;

COMPONENT FILTER_a8237
    PORT (in1 : IN std_logic; y : OUT std_logic);
END COMPONENT;

BEGIN

PROCESS(ain(0), ain(1), ain(2), ain(3), clk, dbin(0), dbin(1), dbin(2), dbin(3),
          dbin(4), dbin(5), dbin(6), dbin(7), dreq(0), dreq(1), dreq(2), dreq(3),
          hlda, ncs, neopin, niorin, niowin, ready, reset)
BEGIN
    ASSERT ain(0) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on ain(0)"
        SEVERITY Warning;
    ASSERT ain(1) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on ain(1)"
        SEVERITY Warning;
    ASSERT ain(2) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on ain(2)"
        SEVERITY Warning;
    ASSERT ain(3) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on ain(3)"
        SEVERITY Warning;
    ASSERT clk /= 'X' OR Now = 0 ns
        REPORT "Unknown value on clk"
        SEVERITY Warning;
    ASSERT dbin(0) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(0)"
        SEVERITY Warning;
    ASSERT dbin(1) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(1)"
        SEVERITY Warning;
    ASSERT dbin(2) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(2)"
        SEVERITY Warning;
    ASSERT dbin(3) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(3)"
        SEVERITY Warning;
    ASSERT dbin(4) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(4)"
        SEVERITY Warning;
    ASSERT dbin(5) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(5)"
        SEVERITY Warning;
    ASSERT dbin(6) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(6)"
        SEVERITY Warning;
    ASSERT dbin(7) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dbin(7)"
        SEVERITY Warning;
    ASSERT dreq(0) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dreq(0)"
        SEVERITY Warning;
    ASSERT dreq(1) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dreq(1)"
        SEVERITY Warning;
    ASSERT dreq(2) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dreq(2)"
        SEVERITY Warning;
    ASSERT dreq(3) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on dreq(3)"
        SEVERITY Warning;
    ASSERT hlda /= 'X' OR Now = 0 ns
        REPORT "Unknown value on hlda"
        SEVERITY Warning;
    ASSERT ncs /= 'X' OR Now = 0 ns
        REPORT "Unknown value on ncs"
        SEVERITY Warning;
    ASSERT neopin /= 'X' OR Now = 0 ns
        REPORT "Unknown value on neopin"
        SEVERITY Warning;
    ASSERT niorin /= 'X' OR Now = 0 ns
        REPORT "Unknown value on niorin"
        SEVERITY Warning;
    ASSERT niowin /= 'X' OR Now = 0 ns
        REPORT "Unknown value on niowin"
        SEVERITY Warning;
    ASSERT ready /= 'X' OR Now = 0 ns
        REPORT "Unknown value on ready"
        SEVERITY Warning;
    ASSERT reset /= 'X' OR Now = 0 ns
        REPORT "Unknown value on reset"
        SEVERITY Warning;
END PROCESS;

tribuf_2: TRIBUF_a8237

    PORT MAP (IN1 => n_153, OE => vcc, Y => dbout(0));
tribuf_4: TRIBUF_a8237

    PORT MAP (IN1 => n_160, OE => vcc, Y => dbout(1));
tribuf_6: TRIBUF_a8237

    PORT MAP (IN1 => n_167, OE => vcc, Y => dbout(2));
tribuf_8: TRIBUF_a8237

    PORT MAP (IN1 => n_174, OE => vcc, Y => dbout(3));
tribuf_10: TRIBUF_a8237

    PORT MAP (IN1 => n_181, OE => vcc, Y => dbout(4));
tribuf_12: TRIBUF_a8237

    PORT MAP (IN1 => n_188, OE => vcc, Y => dbout(5));
tribuf_14: TRIBUF_a8237

    PORT MAP (IN1 => n_195, OE => vcc, Y => dbout(6));
tribuf_16: TRIBUF_a8237

    PORT MAP (IN1 => n_202, OE => vcc, Y => dbout(7));
tribuf_18: TRIBUF_a8237

    PORT MAP (IN1 => n_209, OE => vcc, Y => dack(0));
tribuf_20: TRIBUF_a8237

    PORT MAP (IN1 => n_216, OE => vcc, Y => dack(1));
tribuf_22: TRIBUF_a8237

    PORT MAP (IN1 => n_223, OE => vcc, Y => dack(2));
tribuf_24: TRIBUF_a8237

    PORT MAP (IN1 => n_230, OE => vcc, Y => dack(3));
tribuf_26: TRIBUF_a8237

    PORT MAP (IN1 => n_237, OE => vcc, Y => aout(0));
tribuf_28: TRIBUF_a8237

    PORT MAP (IN1 => n_244, OE => vcc, Y => aout(1));
tribuf_30: TRIBUF_a8237

    PORT MAP (IN1 => n_251, OE => vcc, Y => aout(2));
tribuf_32: TRIBUF_a8237

    PORT MAP (IN1 => n_258, OE => vcc, Y => aout(3));
tribuf_34: TRIBUF_a8237

    PORT MAP (IN1 => n_265, OE => vcc, Y => aout(4));
tribuf_36: TRIBUF_a8237

    PORT MAP (IN1 => n_272, OE => vcc, Y => aout(5));
tribuf_38: TRIBUF_a8237

    PORT MAP (IN1 => n_279, OE => vcc, Y => aout(6));
tribuf_40: TRIBUF_a8237

    PORT MAP (IN1 => n_286, OE => vcc, Y => aout(7));
tribuf_42: TRIBUF_a8237

    PORT MAP (IN1 => n_293, OE => vcc, Y => nmemw);
tribuf_44: TRIBUF_a8237

    PORT MAP (IN1 => n_300, OE => vcc, Y => nmemr);
tribuf_46: TRIBUF_a8237

    PORT MAP (IN1 => n_307, OE => vcc, Y => niowout);
tribuf_48: TRIBUF_a8237

    PORT MAP (IN1 => n_314, OE => vcc, Y => niorout);
tribuf_50: TRIBUF_a8237

    PORT MAP (IN1 => n_321, OE => vcc, Y => neopout);
tribuf_52: TRIBUF_a8237

    PORT MAP (IN1 => n_328, OE => vcc, Y => hrq);
tribuf_54: TRIBUF_a8237

    PORT MAP (IN1 => n_335, OE => vcc, Y => dmaenable);
tribuf_56: TRIBUF_a8237

    PORT MAP (IN1 => n_342, OE => vcc, Y => dben);
tribuf_58: TRIBUF_a8237

    PORT MAP (IN1 => n_349, OE => vcc, Y => aen);
tribuf_60: TRIBUF_a8237

    PORT MAP (IN1 => n_356, OE => vcc, Y => adstb);
delay_61: n_153  <= TRANSPORT n_154  ;
xor2_62: n_154 <=  n_155  XOR n_159;
or1_63: n_155 <=  n_156;
and1_64: n_156 <=  n_157;
delay_65: n_157  <= TRANSPORT a_G956  ;
and1_66: n_159 <=  gnd;
delay_67: n_160  <= TRANSPORT n_161  ;
xor2_68: n_161 <=  n_162  XOR n_166;
or1_69: n_162 <=  n_163;
and1_70: n_163 <=  n_164;
delay_71: n_164  <= TRANSPORT a_G1027  ;
and1_72: n_166 <=  gnd;
delay_73: n_167  <= TRANSPORT n_168  ;
xor2_74: n_168 <=  n_169  XOR n_173;
or1_75: n_169 <=  n_170;
and1_76: n_170 <=  n_171;
delay_77: n_171  <= TRANSPORT a_G200  ;
and1_78: n_173 <=  gnd;
delay_79: n_174  <= TRANSPORT n_175  ;
xor2_80: n_175 <=  n_176  XOR n_180;
or1_81: n_176 <=  n_177;
and1_82: n_177 <=  n_178;
delay_83: n_178  <= TRANSPORT a_G186  ;
and1_84: n_180 <=  gnd;
delay_85: n_181  <= TRANSPORT n_182  ;
xor2_86: n_182 <=  n_183  XOR n_187;
or1_87: n_183 <=  n_184;
and1_88: n_184 <=  n_185;
delay_89: n_185  <= TRANSPORT a_G993  ;
and1_90: n_187 <=  gnd;
delay_91: n_188  <= TRANSPORT n_189  ;
xor2_92: n_189 <=  n_190  XOR n_194;
or1_93: n_190 <=  n_191;
and1_94: n_191 <=  n_192;
delay_95: n_192  <= TRANSPORT a_G917  ;
and1_96: n_194 <=  gnd;
delay_97: n_195  <= TRANSPORT n_196  ;
xor2_98: n_196 <=  n_197  XOR n_201;
or1_99: n_197 <=  n_198;
and1_100: n_198 <=  n_199;
delay_101: n_199  <= TRANSPORT a_G142  ;
and1_102: n_201 <=  gnd;
delay_103: n_202  <= TRANSPORT n_203  ;
xor2_104: n_203 <=  n_204  XOR n_208;
or1_105: n_204 <=  n_205;
and1_106: n_205 <=  n_206;
delay_107: n_206  <= TRANSPORT a_G1389  ;
and1_108: n_208 <=  gnd;
delay_109: n_209  <= TRANSPORT n_210  ;
xor2_110: n_210 <=  n_211  XOR n_215;
or1_111: n_211 <=  n_212;
and1_112: n_212 <=  n_213;
delay_113: n_213  <= TRANSPORT a_G503  ;
and1_114: n_215 <=  gnd;
delay_115: n_216  <= TRANSPORT n_217  ;
xor2_116: n_217 <=  n_218  XOR n_222;
or1_117: n_218 <=  n_219;
and1_118: n_219 <=  n_220;
delay_119: n_220  <= TRANSPORT a_G502  ;
and1_120: n_222 <=  gnd;
delay_121: n_223  <= TRANSPORT n_224  ;
xor2_122: n_224 <=  n_225  XOR n_229;
or1_123: n_225 <=  n_226;
and1_124: n_226 <=  n_227;
delay_125: n_227  <= TRANSPORT a_G1464  ;
and1_126: n_229 <=  gnd;
delay_127: n_230  <= TRANSPORT n_231  ;
xor2_128: n_231 <=  n_232  XOR n_236;
or1_129: n_232 <=  n_233;
and1_130: n_233 <=  n_234;
delay_131: n_234  <= TRANSPORT a_G1463  ;
and1_132: n_236 <=  gnd;
delay_133: n_237  <= TRANSPORT n_238  ;
xor2_134: n_238 <=  n_239  XOR n_243;
or1_135: n_239 <=  n_240;
and1_136: n_240 <=  n_241;
delay_137: n_241  <= TRANSPORT a_LC7_D18  ;
and1_138: n_243 <=  gnd;
delay_139: n_244  <= TRANSPORT n_245  ;
xor2_140: n_245 <=  n_246  XOR n_250;
or1_141: n_246 <=  n_247;
and1_142: n_247 <=  n_248;
delay_143: n_248  <= TRANSPORT a_LC7_C17  ;
and1_144: n_250 <=  gnd;
delay_145: n_251  <= TRANSPORT n_252  ;
xor2_146: n_252 <=  n_253  XOR n_257;
or1_147: n_253 <=  n_254;
and1_148: n_254 <=  n_255;
delay_149: n_255  <= TRANSPORT a_LC4_C16  ;
and1_150: n_257 <=  gnd;
delay_151: n_258  <= TRANSPORT n_259  ;
xor2_152: n_259 <=  n_260  XOR n_264;
or1_153: n_260 <=  n_261;
and1_154: n_261 <=  n_262;
delay_155: n_262  <= TRANSPORT a_LC2_C24  ;
and1_156: n_264 <=  gnd;
delay_157: n_265  <= TRANSPORT n_266  ;
xor2_158: n_266 <=  n_267  XOR n_271;
or1_159: n_267 <=  n_268;
and1_160: n_268 <=  n_269;
delay_161: n_269  <= TRANSPORT a_LC1_C16  ;
and1_162: n_271 <=  gnd;
delay_163: n_272  <= TRANSPORT n_273  ;
xor2_164: n_273 <=  n_274  XOR n_278;
or1_165: n_274 <=  n_275;
and1_166: n_275 <=  n_276;
delay_167: n_276  <= TRANSPORT a_LC3_F6  ;
and1_168: n_278 <=  gnd;
delay_169: n_279  <= TRANSPORT n_280  ;
xor2_170: n_280 <=  n_281  XOR n_285;
or1_171: n_281 <=  n_282;
and1_172: n_282 <=  n_283;
delay_173: n_283  <= TRANSPORT a_LC4_F10  ;
and1_174: n_285 <=  gnd;
delay_175: n_286  <= TRANSPORT n_287  ;
xor2_176: n_287 <=  n_288  XOR n_292;
or1_177: n_288 <=  n_289;
and1_178: n_289 <=  n_290;
delay_179: n_290  <= TRANSPORT a_LC5_D27  ;
and1_180: n_292 <=  gnd;
delay_181: n_293  <= TRANSPORT n_294  ;
xor2_182: n_294 <=  n_295  XOR n_299;
or1_183: n_295 <=  n_296;
and1_184: n_296 <=  n_297;
delay_185: n_297  <= TRANSPORT a_SNMEMW  ;
and1_186: n_299 <=  gnd;
delay_187: n_300  <= TRANSPORT n_301  ;
xor2_188: n_301 <=  n_302  XOR n_306;
or1_189: n_302 <=  n_303;
and1_190: n_303 <=  n_304;
inv_191: n_304  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
and1_192: n_306 <=  gnd;
delay_193: n_307  <= TRANSPORT n_308  ;
xor2_194: n_308 <=  n_309  XOR n_313;
or1_195: n_309 <=  n_310;
and1_196: n_310 <=  n_311;
delay_197: n_311  <= TRANSPORT a_SNIOWOUT  ;
and1_198: n_313 <=  gnd;
delay_199: n_314  <= TRANSPORT n_315  ;
xor2_200: n_315 <=  n_316  XOR n_320;
or1_201: n_316 <=  n_317;
and1_202: n_317 <=  n_318;
delay_203: n_318  <= TRANSPORT a_SNIOROUT  ;
and1_204: n_320 <=  gnd;
delay_205: n_321  <= TRANSPORT n_322  ;
xor2_206: n_322 <=  n_323  XOR n_327;
or1_207: n_323 <=  n_324;
and1_208: n_324 <=  n_325;
inv_209: n_325  <= TRANSPORT NOT a_SNEOPOUT_aNOT  ;
and1_210: n_327 <=  gnd;
delay_211: n_328  <= TRANSPORT n_329  ;
xor2_212: n_329 <=  n_330  XOR n_334;
or1_213: n_330 <=  n_331;
and1_214: n_331 <=  n_332;
delay_215: n_332  <= TRANSPORT a_SHRQ  ;
and1_216: n_334 <=  gnd;
delay_217: n_335  <= TRANSPORT n_336  ;
xor2_218: n_336 <=  n_337  XOR n_341;
or1_219: n_337 <=  n_338;
and1_220: n_338 <=  n_339;
inv_221: n_339  <= TRANSPORT NOT a_SAEN_aNOT  ;
and1_222: n_341 <=  gnd;
delay_223: n_342  <= TRANSPORT n_343  ;
xor2_224: n_343 <=  n_344  XOR n_348;
or1_225: n_344 <=  n_345;
and1_226: n_345 <=  n_346;
delay_227: n_346  <= TRANSPORT a_SDBEN  ;
and1_228: n_348 <=  gnd;
delay_229: n_349  <= TRANSPORT n_350  ;
xor2_230: n_350 <=  n_351  XOR n_355;
or1_231: n_351 <=  n_352;
and1_232: n_352 <=  n_353;
inv_233: n_353  <= TRANSPORT NOT a_LC6_B16_aNOT  ;
and1_234: n_355 <=  gnd;
delay_235: n_356  <= TRANSPORT n_357  ;
xor2_236: n_357 <=  n_358  XOR n_362;
or1_237: n_358 <=  n_359;
and1_238: n_359 <=  n_360;
delay_239: n_360  <= TRANSPORT a_SADSTB  ;
and1_240: n_362 <=  gnd;
dff_241: DFF_a8237

    PORT MAP ( D => a_EQ1030, CLK => a_SCH2BWORDOUT_F3_G_aCLK, CLRN => a_SCH2BWORDOUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F3_G);
inv_242: a_SCH2BWORDOUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_243: a_EQ1030 <=  n_371  XOR n_380;
or2_244: n_371 <=  n_372  OR n_377;
and2_245: n_372 <=  n_373  AND n_375;
inv_246: n_373  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_247: n_375  <= TRANSPORT dbin(3)  ;
and2_248: n_377 <=  n_378  AND n_379;
delay_249: n_378  <= TRANSPORT a_N2574_aNOT  ;
delay_250: n_379  <= TRANSPORT a_SCH2BWORDOUT_F3_G  ;
and1_251: n_380 <=  gnd;
delay_252: n_381  <= TRANSPORT clk  ;
filter_253: FILTER_a8237

    PORT MAP (IN1 => n_381, Y => a_SCH2BWORDOUT_F3_G_aCLK);
dff_254: DFF_a8237

    PORT MAP ( D => a_EQ903, CLK => a_SCH0BWORDOUT_F4_G_aCLK, CLRN => a_SCH0BWORDOUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F4_G);
inv_255: a_SCH0BWORDOUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_256: a_EQ903 <=  n_391  XOR n_400;
or2_257: n_391 <=  n_392  OR n_397;
and2_258: n_392 <=  n_393  AND n_395;
inv_259: n_393  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_260: n_395  <= TRANSPORT dbin(4)  ;
and2_261: n_397 <=  n_398  AND n_399;
delay_262: n_398  <= TRANSPORT a_N2578_aNOT  ;
delay_263: n_399  <= TRANSPORT a_SCH0BWORDOUT_F4_G  ;
and1_264: n_400 <=  gnd;
delay_265: n_401  <= TRANSPORT clk  ;
filter_266: FILTER_a8237

    PORT MAP (IN1 => n_401, Y => a_SCH0BWORDOUT_F4_G_aCLK);
dff_267: DFF_a8237

    PORT MAP ( D => a_EQ1095, CLK => a_SCH3BWORDOUT_F4_G_aCLK, CLRN => a_SCH3BWORDOUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F4_G);
inv_268: a_SCH3BWORDOUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_269: a_EQ1095 <=  n_410  XOR n_418;
or2_270: n_410 <=  n_411  OR n_415;
and2_271: n_411 <=  n_412  AND n_414;
inv_272: n_412  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_273: n_414  <= TRANSPORT dbin(4)  ;
and2_274: n_415 <=  n_416  AND n_417;
delay_275: n_416  <= TRANSPORT a_N2572_aNOT  ;
delay_276: n_417  <= TRANSPORT a_SCH3BWORDOUT_F4_G  ;
and1_277: n_418 <=  gnd;
delay_278: n_419  <= TRANSPORT clk  ;
filter_279: FILTER_a8237

    PORT MAP (IN1 => n_419, Y => a_SCH3BWORDOUT_F4_G_aCLK);
dff_280: DFF_a8237

    PORT MAP ( D => a_EQ1031, CLK => a_SCH2BWORDOUT_F4_G_aCLK, CLRN => a_SCH2BWORDOUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F4_G);
inv_281: a_SCH2BWORDOUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_282: a_EQ1031 <=  n_428  XOR n_435;
or2_283: n_428 <=  n_429  OR n_432;
and2_284: n_429 <=  n_430  AND n_431;
inv_285: n_430  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_286: n_431  <= TRANSPORT dbin(4)  ;
and2_287: n_432 <=  n_433  AND n_434;
delay_288: n_433  <= TRANSPORT a_N2574_aNOT  ;
delay_289: n_434  <= TRANSPORT a_SCH2BWORDOUT_F4_G  ;
and1_290: n_435 <=  gnd;
delay_291: n_436  <= TRANSPORT clk  ;
filter_292: FILTER_a8237

    PORT MAP (IN1 => n_436, Y => a_SCH2BWORDOUT_F4_G_aCLK);
dff_293: DFF_a8237

    PORT MAP ( D => a_EQ967, CLK => a_SCH1BWORDOUT_F4_G_aCLK, CLRN => a_SCH1BWORDOUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F4_G);
inv_294: a_SCH1BWORDOUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_295: a_EQ967 <=  n_445  XOR n_453;
or2_296: n_445 <=  n_446  OR n_450;
and2_297: n_446 <=  n_447  AND n_449;
inv_298: n_447  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_299: n_449  <= TRANSPORT dbin(4)  ;
and2_300: n_450 <=  n_451  AND n_452;
delay_301: n_451  <= TRANSPORT a_N2576_aNOT  ;
delay_302: n_452  <= TRANSPORT a_SCH1BWORDOUT_F4_G  ;
and1_303: n_453 <=  gnd;
delay_304: n_454  <= TRANSPORT clk  ;
filter_305: FILTER_a8237

    PORT MAP (IN1 => n_454, Y => a_SCH1BWORDOUT_F4_G_aCLK);
delay_306: a_N2352  <= TRANSPORT a_EQ556  ;
xor2_307: a_EQ556 <=  n_458  XOR n_471;
or4_308: n_458 <=  n_459  OR n_462  OR n_465  OR n_468;
and1_309: n_459 <=  n_460;
delay_310: n_460  <= TRANSPORT ain(2)  ;
and1_311: n_462 <=  n_463;
inv_312: n_463  <= TRANSPORT NOT ain(1)  ;
and1_313: n_465 <=  n_466;
delay_314: n_466  <= TRANSPORT ain(0)  ;
and1_315: n_468 <=  n_469;
delay_316: n_469  <= TRANSPORT ain(3)  ;
and1_317: n_471 <=  gnd;
delay_318: a_N2585_aNOT  <= TRANSPORT a_EQ638  ;
xor2_319: a_EQ638 <=  n_474  XOR n_480;
or2_320: n_474 <=  n_475  OR n_477;
and1_321: n_475 <=  n_476;
delay_322: n_476  <= TRANSPORT a_N2352  ;
and1_323: n_477 <=  n_478;
delay_324: n_478  <= TRANSPORT a_LC3_D22  ;
and1_325: n_480 <=  gnd;
dff_326: DFF_a8237

    PORT MAP ( D => a_EQ959, CLK => a_SCH1BAROUT_F12_G_aCLK, CLRN => a_SCH1BAROUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F12_G);
inv_327: a_SCH1BAROUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_328: a_EQ959 <=  n_488  XOR n_495;
or2_329: n_488 <=  n_489  OR n_492;
and2_330: n_489 <=  n_490  AND n_491;
inv_331: n_490  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_332: n_491  <= TRANSPORT dbin(4)  ;
and2_333: n_492 <=  n_493  AND n_494;
delay_334: n_493  <= TRANSPORT a_N2585_aNOT  ;
delay_335: n_494  <= TRANSPORT a_SCH1BAROUT_F12_G  ;
and1_336: n_495 <=  gnd;
delay_337: n_496  <= TRANSPORT clk  ;
filter_338: FILTER_a8237

    PORT MAP (IN1 => n_496, Y => a_SCH1BAROUT_F12_G_aCLK);
dff_339: DFF_a8237

    PORT MAP ( D => a_EQ960, CLK => a_SCH1BAROUT_F13_G_aCLK, CLRN => a_SCH1BAROUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F13_G);
inv_340: a_SCH1BAROUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_341: a_EQ960 <=  n_505  XOR n_513;
or2_342: n_505 <=  n_506  OR n_510;
and2_343: n_506 <=  n_507  AND n_508;
inv_344: n_507  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_345: n_508  <= TRANSPORT dbin(5)  ;
and2_346: n_510 <=  n_511  AND n_512;
delay_347: n_511  <= TRANSPORT a_N2585_aNOT  ;
delay_348: n_512  <= TRANSPORT a_SCH1BAROUT_F13_G  ;
and1_349: n_513 <=  gnd;
delay_350: n_514  <= TRANSPORT clk  ;
filter_351: FILTER_a8237

    PORT MAP (IN1 => n_514, Y => a_SCH1BAROUT_F13_G_aCLK);
dff_352: DFF_a8237

    PORT MAP ( D => a_EQ1033, CLK => a_SCH2BWORDOUT_F6_G_aCLK, CLRN => a_SCH2BWORDOUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F6_G);
inv_353: a_SCH2BWORDOUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_354: a_EQ1033 <=  n_523  XOR n_531;
or2_355: n_523 <=  n_524  OR n_528;
and2_356: n_524 <=  n_525  AND n_526;
inv_357: n_525  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_358: n_526  <= TRANSPORT dbin(6)  ;
and2_359: n_528 <=  n_529  AND n_530;
delay_360: n_529  <= TRANSPORT a_N2574_aNOT  ;
delay_361: n_530  <= TRANSPORT a_SCH2BWORDOUT_F6_G  ;
and1_362: n_531 <=  gnd;
delay_363: n_532  <= TRANSPORT clk  ;
filter_364: FILTER_a8237

    PORT MAP (IN1 => n_532, Y => a_SCH2BWORDOUT_F6_G_aCLK);
dff_365: DFF_a8237

    PORT MAP ( D => a_EQ969, CLK => a_SCH1BWORDOUT_F6_G_aCLK, CLRN => a_SCH1BWORDOUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F6_G);
inv_366: a_SCH1BWORDOUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_367: a_EQ969 <=  n_541  XOR n_548;
or2_368: n_541 <=  n_542  OR n_545;
and2_369: n_542 <=  n_543  AND n_544;
inv_370: n_543  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_371: n_544  <= TRANSPORT dbin(6)  ;
and2_372: n_545 <=  n_546  AND n_547;
delay_373: n_546  <= TRANSPORT a_N2576_aNOT  ;
delay_374: n_547  <= TRANSPORT a_SCH1BWORDOUT_F6_G  ;
and1_375: n_548 <=  gnd;
delay_376: n_549  <= TRANSPORT clk  ;
filter_377: FILTER_a8237

    PORT MAP (IN1 => n_549, Y => a_SCH1BWORDOUT_F6_G_aCLK);
dff_378: DFF_a8237

    PORT MAP ( D => a_EQ905, CLK => a_SCH0BWORDOUT_F6_G_aCLK, CLRN => a_SCH0BWORDOUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F6_G);
inv_379: a_SCH0BWORDOUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_380: a_EQ905 <=  n_558  XOR n_565;
or2_381: n_558 <=  n_559  OR n_562;
and2_382: n_559 <=  n_560  AND n_561;
inv_383: n_560  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_384: n_561  <= TRANSPORT dbin(6)  ;
and2_385: n_562 <=  n_563  AND n_564;
delay_386: n_563  <= TRANSPORT a_N2578_aNOT  ;
delay_387: n_564  <= TRANSPORT a_SCH0BWORDOUT_F6_G  ;
and1_388: n_565 <=  gnd;
delay_389: n_566  <= TRANSPORT clk  ;
filter_390: FILTER_a8237

    PORT MAP (IN1 => n_566, Y => a_SCH0BWORDOUT_F6_G_aCLK);
delay_391: a_N77_aNOT  <= TRANSPORT a_EQ194  ;
xor2_392: a_EQ194 <=  n_570  XOR n_579;
or4_393: n_570 <=  n_571  OR n_573  OR n_575  OR n_577;
and1_394: n_571 <=  n_572;
delay_395: n_572  <= TRANSPORT ain(0)  ;
and1_396: n_573 <=  n_574;
delay_397: n_574  <= TRANSPORT ain(3)  ;
and1_398: n_575 <=  n_576;
inv_399: n_576  <= TRANSPORT NOT ain(2)  ;
and1_400: n_577 <=  n_578;
delay_401: n_578  <= TRANSPORT ain(1)  ;
and1_402: n_579 <=  gnd;
delay_403: a_N2583_aNOT  <= TRANSPORT a_EQ636  ;
xor2_404: a_EQ636 <=  n_582  XOR n_587;
or2_405: n_582 <=  n_583  OR n_585;
and1_406: n_583 <=  n_584;
delay_407: n_584  <= TRANSPORT a_N77_aNOT  ;
and1_408: n_585 <=  n_586;
delay_409: n_586  <= TRANSPORT a_LC3_D22  ;
and1_410: n_587 <=  gnd;
dff_411: DFF_a8237

    PORT MAP ( D => a_EQ1025, CLK => a_SCH2BAROUT_F14_G_aCLK, CLRN => a_SCH2BAROUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F14_G);
inv_412: a_SCH2BAROUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_413: a_EQ1025 <=  n_595  XOR n_602;
or2_414: n_595 <=  n_596  OR n_599;
and2_415: n_596 <=  n_597  AND n_598;
inv_416: n_597  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_417: n_598  <= TRANSPORT dbin(6)  ;
and2_418: n_599 <=  n_600  AND n_601;
delay_419: n_600  <= TRANSPORT a_N2583_aNOT  ;
delay_420: n_601  <= TRANSPORT a_SCH2BAROUT_F14_G  ;
and1_421: n_602 <=  gnd;
delay_422: n_603  <= TRANSPORT clk  ;
filter_423: FILTER_a8237

    PORT MAP (IN1 => n_603, Y => a_SCH2BAROUT_F14_G_aCLK);
dff_424: DFF_a8237

    PORT MAP ( D => a_EQ961, CLK => a_SCH1BAROUT_F14_G_aCLK, CLRN => a_SCH1BAROUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F14_G);
inv_425: a_SCH1BAROUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_426: a_EQ961 <=  n_612  XOR n_619;
or2_427: n_612 <=  n_613  OR n_616;
and2_428: n_613 <=  n_614  AND n_615;
inv_429: n_614  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_430: n_615  <= TRANSPORT dbin(6)  ;
and2_431: n_616 <=  n_617  AND n_618;
delay_432: n_617  <= TRANSPORT a_N2585_aNOT  ;
delay_433: n_618  <= TRANSPORT a_SCH1BAROUT_F14_G  ;
and1_434: n_619 <=  gnd;
delay_435: n_620  <= TRANSPORT clk  ;
filter_436: FILTER_a8237

    PORT MAP (IN1 => n_620, Y => a_SCH1BAROUT_F14_G_aCLK);
dff_437: DFF_a8237

    PORT MAP ( D => a_EQ970, CLK => a_SCH1BWORDOUT_F7_G_aCLK, CLRN => a_SCH1BWORDOUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F7_G);
inv_438: a_SCH1BWORDOUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_439: a_EQ970 <=  n_629  XOR n_637;
or2_440: n_629 <=  n_630  OR n_634;
and2_441: n_630 <=  n_631  AND n_632;
inv_442: n_631  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_443: n_632  <= TRANSPORT dbin(7)  ;
and2_444: n_634 <=  n_635  AND n_636;
delay_445: n_635  <= TRANSPORT a_N2576_aNOT  ;
delay_446: n_636  <= TRANSPORT a_SCH1BWORDOUT_F7_G  ;
and1_447: n_637 <=  gnd;
delay_448: n_638  <= TRANSPORT clk  ;
filter_449: FILTER_a8237

    PORT MAP (IN1 => n_638, Y => a_SCH1BWORDOUT_F7_G_aCLK);
delay_450: a_N2573_aNOT  <= TRANSPORT a_EQ626  ;
xor2_451: a_EQ626 <=  n_642  XOR n_652;
or3_452: n_642 <=  n_643  OR n_646  OR n_649;
and1_453: n_643 <=  n_644;
inv_454: n_644  <= TRANSPORT NOT bytepointer  ;
and1_455: n_646 <=  n_647;
delay_456: n_647  <= TRANSPORT a_N87  ;
and1_457: n_649 <=  n_650;
delay_458: n_650  <= TRANSPORT a_N2347  ;
and1_459: n_652 <=  gnd;
dff_460: DFF_a8237

    PORT MAP ( D => a_EQ1102, CLK => a_SCH3BWORDOUT_F11_G_aCLK, CLRN => a_SCH3BWORDOUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F11_G);
inv_461: a_SCH3BWORDOUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_462: a_EQ1102 <=  n_660  XOR n_667;
or2_463: n_660 <=  n_661  OR n_664;
and2_464: n_661 <=  n_662  AND n_663;
inv_465: n_662  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_466: n_663  <= TRANSPORT dbin(3)  ;
and2_467: n_664 <=  n_665  AND n_666;
delay_468: n_665  <= TRANSPORT a_N2573_aNOT  ;
delay_469: n_666  <= TRANSPORT a_SCH3BWORDOUT_F11_G  ;
and1_470: n_667 <=  gnd;
delay_471: n_668  <= TRANSPORT clk  ;
filter_472: FILTER_a8237

    PORT MAP (IN1 => n_668, Y => a_SCH3BWORDOUT_F11_G_aCLK);
dff_473: DFF_a8237

    PORT MAP ( D => a_EQ974, CLK => a_SCH1BWORDOUT_F11_G_aCLK, CLRN => a_SCH1BWORDOUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F11_G);
inv_474: a_SCH1BWORDOUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_475: a_EQ974 <=  n_677  XOR n_685;
or2_476: n_677 <=  n_678  OR n_682;
and2_477: n_678 <=  n_679  AND n_681;
inv_478: n_679  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_479: n_681  <= TRANSPORT dbin(3)  ;
and2_480: n_682 <=  n_683  AND n_684;
delay_481: n_683  <= TRANSPORT a_N2577_aNOT  ;
delay_482: n_684  <= TRANSPORT a_SCH1BWORDOUT_F11_G  ;
and1_483: n_685 <=  gnd;
delay_484: n_686  <= TRANSPORT clk  ;
filter_485: FILTER_a8237

    PORT MAP (IN1 => n_686, Y => a_SCH1BWORDOUT_F11_G_aCLK);
dff_486: DFF_a8237

    PORT MAP ( D => a_EQ1038, CLK => a_SCH2BWORDOUT_F11_G_aCLK, CLRN => a_SCH2BWORDOUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F11_G);
inv_487: a_SCH2BWORDOUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_488: a_EQ1038 <=  n_695  XOR n_707;
or3_489: n_695 <=  n_696  OR n_701  OR n_704;
and3_490: n_696 <=  n_697  AND n_698  AND n_700;
inv_491: n_697  <= TRANSPORT NOT a_LC3_D22  ;
inv_492: n_698  <= TRANSPORT NOT a_N62_aNOT  ;
delay_493: n_700  <= TRANSPORT dbin(3)  ;
and2_494: n_701 <=  n_702  AND n_703;
delay_495: n_702  <= TRANSPORT a_N62_aNOT  ;
delay_496: n_703  <= TRANSPORT a_SCH2BWORDOUT_F11_G  ;
and2_497: n_704 <=  n_705  AND n_706;
delay_498: n_705  <= TRANSPORT a_LC3_D22  ;
delay_499: n_706  <= TRANSPORT a_SCH2BWORDOUT_F11_G  ;
and1_500: n_707 <=  gnd;
delay_501: n_708  <= TRANSPORT clk  ;
filter_502: FILTER_a8237

    PORT MAP (IN1 => n_708, Y => a_SCH2BWORDOUT_F11_G_aCLK);
dff_503: DFF_a8237

    PORT MAP ( D => a_EQ910, CLK => a_SCH0BWORDOUT_F11_G_aCLK, CLRN => a_SCH0BWORDOUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F11_G);
inv_504: a_SCH0BWORDOUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_505: a_EQ910 <=  n_717  XOR n_729;
or3_506: n_717 <=  n_718  OR n_723  OR n_726;
and3_507: n_718 <=  n_719  AND n_720  AND n_722;
inv_508: n_719  <= TRANSPORT NOT a_LC3_D22  ;
inv_509: n_720  <= TRANSPORT NOT a_N2353  ;
delay_510: n_722  <= TRANSPORT dbin(3)  ;
and2_511: n_723 <=  n_724  AND n_725;
delay_512: n_724  <= TRANSPORT a_N2353  ;
delay_513: n_725  <= TRANSPORT a_SCH0BWORDOUT_F11_G  ;
and2_514: n_726 <=  n_727  AND n_728;
delay_515: n_727  <= TRANSPORT a_LC3_D22  ;
delay_516: n_728  <= TRANSPORT a_SCH0BWORDOUT_F11_G  ;
and1_517: n_729 <=  gnd;
delay_518: n_730  <= TRANSPORT clk  ;
filter_519: FILTER_a8237

    PORT MAP (IN1 => n_730, Y => a_SCH0BWORDOUT_F11_G_aCLK);
dff_520: DFF_a8237

    PORT MAP ( D => a_EQ1103, CLK => a_SCH3BWORDOUT_F12_G_aCLK, CLRN => a_SCH3BWORDOUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F12_G);
inv_521: a_SCH3BWORDOUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_522: a_EQ1103 <=  n_739  XOR n_746;
or2_523: n_739 <=  n_740  OR n_743;
and2_524: n_740 <=  n_741  AND n_742;
inv_525: n_741  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_526: n_742  <= TRANSPORT dbin(4)  ;
and2_527: n_743 <=  n_744  AND n_745;
delay_528: n_744  <= TRANSPORT a_N2573_aNOT  ;
delay_529: n_745  <= TRANSPORT a_SCH3BWORDOUT_F12_G  ;
and1_530: n_746 <=  gnd;
delay_531: n_747  <= TRANSPORT clk  ;
filter_532: FILTER_a8237

    PORT MAP (IN1 => n_747, Y => a_SCH3BWORDOUT_F12_G_aCLK);
dff_533: DFF_a8237

    PORT MAP ( D => a_EQ911, CLK => a_SCH0BWORDOUT_F12_G_aCLK, CLRN => a_SCH0BWORDOUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F12_G);
inv_534: a_SCH0BWORDOUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_535: a_EQ911 <=  n_756  XOR n_767;
or3_536: n_756 <=  n_757  OR n_761  OR n_764;
and3_537: n_757 <=  n_758  AND n_759  AND n_760;
inv_538: n_758  <= TRANSPORT NOT a_LC3_D22  ;
inv_539: n_759  <= TRANSPORT NOT a_N2353  ;
delay_540: n_760  <= TRANSPORT dbin(4)  ;
and2_541: n_761 <=  n_762  AND n_763;
delay_542: n_762  <= TRANSPORT a_N2353  ;
delay_543: n_763  <= TRANSPORT a_SCH0BWORDOUT_F12_G  ;
and2_544: n_764 <=  n_765  AND n_766;
delay_545: n_765  <= TRANSPORT a_LC3_D22  ;
delay_546: n_766  <= TRANSPORT a_SCH0BWORDOUT_F12_G  ;
and1_547: n_767 <=  gnd;
delay_548: n_768  <= TRANSPORT clk  ;
filter_549: FILTER_a8237

    PORT MAP (IN1 => n_768, Y => a_SCH0BWORDOUT_F12_G_aCLK);
dff_550: DFF_a8237

    PORT MAP ( D => a_EQ1039, CLK => a_SCH2BWORDOUT_F12_G_aCLK, CLRN => a_SCH2BWORDOUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F12_G);
inv_551: a_SCH2BWORDOUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_552: a_EQ1039 <=  n_777  XOR n_788;
or3_553: n_777 <=  n_778  OR n_782  OR n_785;
and3_554: n_778 <=  n_779  AND n_780  AND n_781;
inv_555: n_779  <= TRANSPORT NOT a_LC3_D22  ;
inv_556: n_780  <= TRANSPORT NOT a_N62_aNOT  ;
delay_557: n_781  <= TRANSPORT dbin(4)  ;
and2_558: n_782 <=  n_783  AND n_784;
delay_559: n_783  <= TRANSPORT a_N62_aNOT  ;
delay_560: n_784  <= TRANSPORT a_SCH2BWORDOUT_F12_G  ;
and2_561: n_785 <=  n_786  AND n_787;
delay_562: n_786  <= TRANSPORT a_LC3_D22  ;
delay_563: n_787  <= TRANSPORT a_SCH2BWORDOUT_F12_G  ;
and1_564: n_788 <=  gnd;
delay_565: n_789  <= TRANSPORT clk  ;
filter_566: FILTER_a8237

    PORT MAP (IN1 => n_789, Y => a_SCH2BWORDOUT_F12_G_aCLK);
dff_567: DFF_a8237

    PORT MAP ( D => a_EQ975, CLK => a_SCH1BWORDOUT_F12_G_aCLK, CLRN => a_SCH1BWORDOUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F12_G);
inv_568: a_SCH1BWORDOUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_569: a_EQ975 <=  n_798  XOR n_805;
or2_570: n_798 <=  n_799  OR n_802;
and2_571: n_799 <=  n_800  AND n_801;
inv_572: n_800  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_573: n_801  <= TRANSPORT dbin(4)  ;
and2_574: n_802 <=  n_803  AND n_804;
delay_575: n_803  <= TRANSPORT a_N2577_aNOT  ;
delay_576: n_804  <= TRANSPORT a_SCH1BWORDOUT_F12_G  ;
and1_577: n_805 <=  gnd;
delay_578: n_806  <= TRANSPORT clk  ;
filter_579: FILTER_a8237

    PORT MAP (IN1 => n_806, Y => a_SCH1BWORDOUT_F12_G_aCLK);
dff_580: DFF_a8237

    PORT MAP ( D => a_EQ1093, CLK => a_SCH3BWORDOUT_F2_G_aCLK, CLRN => a_SCH3BWORDOUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F2_G);
inv_581: a_SCH3BWORDOUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_582: a_EQ1093 <=  n_815  XOR n_823;
or2_583: n_815 <=  n_816  OR n_820;
and2_584: n_816 <=  n_817  AND n_818;
inv_585: n_817  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_586: n_818  <= TRANSPORT dbin(2)  ;
and2_587: n_820 <=  n_821  AND n_822;
delay_588: n_821  <= TRANSPORT a_N2572_aNOT  ;
delay_589: n_822  <= TRANSPORT a_SCH3BWORDOUT_F2_G  ;
and1_590: n_823 <=  gnd;
delay_591: n_824  <= TRANSPORT clk  ;
filter_592: FILTER_a8237

    PORT MAP (IN1 => n_824, Y => a_SCH3BWORDOUT_F2_G_aCLK);
dff_593: DFF_a8237

    PORT MAP ( D => a_EQ1029, CLK => a_SCH2BWORDOUT_F2_G_aCLK, CLRN => a_SCH2BWORDOUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F2_G);
inv_594: a_SCH2BWORDOUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_595: a_EQ1029 <=  n_833  XOR n_840;
or2_596: n_833 <=  n_834  OR n_837;
and2_597: n_834 <=  n_835  AND n_836;
inv_598: n_835  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_599: n_836  <= TRANSPORT dbin(2)  ;
and2_600: n_837 <=  n_838  AND n_839;
delay_601: n_838  <= TRANSPORT a_N2574_aNOT  ;
delay_602: n_839  <= TRANSPORT a_SCH2BWORDOUT_F2_G  ;
and1_603: n_840 <=  gnd;
delay_604: n_841  <= TRANSPORT clk  ;
filter_605: FILTER_a8237

    PORT MAP (IN1 => n_841, Y => a_SCH2BWORDOUT_F2_G_aCLK);
dff_606: DFF_a8237

    PORT MAP ( D => a_EQ1105, CLK => a_SCH3BWORDOUT_F14_G_aCLK, CLRN => a_SCH3BWORDOUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F14_G);
inv_607: a_SCH3BWORDOUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_608: a_EQ1105 <=  n_850  XOR n_857;
or2_609: n_850 <=  n_851  OR n_854;
and2_610: n_851 <=  n_852  AND n_853;
inv_611: n_852  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_612: n_853  <= TRANSPORT dbin(6)  ;
and2_613: n_854 <=  n_855  AND n_856;
delay_614: n_855  <= TRANSPORT a_N2573_aNOT  ;
delay_615: n_856  <= TRANSPORT a_SCH3BWORDOUT_F14_G  ;
and1_616: n_857 <=  gnd;
delay_617: n_858  <= TRANSPORT clk  ;
filter_618: FILTER_a8237

    PORT MAP (IN1 => n_858, Y => a_SCH3BWORDOUT_F14_G_aCLK);
dff_619: DFF_a8237

    PORT MAP ( D => a_EQ977, CLK => a_SCH1BWORDOUT_F14_G_aCLK, CLRN => a_SCH1BWORDOUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F14_G);
inv_620: a_SCH1BWORDOUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_621: a_EQ977 <=  n_867  XOR n_874;
or2_622: n_867 <=  n_868  OR n_871;
and2_623: n_868 <=  n_869  AND n_870;
inv_624: n_869  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_625: n_870  <= TRANSPORT dbin(6)  ;
and2_626: n_871 <=  n_872  AND n_873;
delay_627: n_872  <= TRANSPORT a_N2577_aNOT  ;
delay_628: n_873  <= TRANSPORT a_SCH1BWORDOUT_F14_G  ;
and1_629: n_874 <=  gnd;
delay_630: n_875  <= TRANSPORT clk  ;
filter_631: FILTER_a8237

    PORT MAP (IN1 => n_875, Y => a_SCH1BWORDOUT_F14_G_aCLK);
dff_632: DFF_a8237

    PORT MAP ( D => a_EQ1041, CLK => a_SCH2BWORDOUT_F14_G_aCLK, CLRN => a_SCH2BWORDOUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F14_G);
inv_633: a_SCH2BWORDOUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_634: a_EQ1041 <=  n_884  XOR n_895;
or3_635: n_884 <=  n_885  OR n_889  OR n_892;
and3_636: n_885 <=  n_886  AND n_887  AND n_888;
inv_637: n_886  <= TRANSPORT NOT a_LC3_D22  ;
inv_638: n_887  <= TRANSPORT NOT a_N62_aNOT  ;
delay_639: n_888  <= TRANSPORT dbin(6)  ;
and2_640: n_889 <=  n_890  AND n_891;
delay_641: n_890  <= TRANSPORT a_N62_aNOT  ;
delay_642: n_891  <= TRANSPORT a_SCH2BWORDOUT_F14_G  ;
and2_643: n_892 <=  n_893  AND n_894;
delay_644: n_893  <= TRANSPORT a_LC3_D22  ;
delay_645: n_894  <= TRANSPORT a_SCH2BWORDOUT_F14_G  ;
and1_646: n_895 <=  gnd;
delay_647: n_896  <= TRANSPORT clk  ;
filter_648: FILTER_a8237

    PORT MAP (IN1 => n_896, Y => a_SCH2BWORDOUT_F14_G_aCLK);
dff_649: DFF_a8237

    PORT MAP ( D => a_EQ913, CLK => a_SCH0BWORDOUT_F14_G_aCLK, CLRN => a_SCH0BWORDOUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F14_G);
inv_650: a_SCH0BWORDOUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_651: a_EQ913 <=  n_905  XOR n_916;
or3_652: n_905 <=  n_906  OR n_910  OR n_913;
and3_653: n_906 <=  n_907  AND n_908  AND n_909;
inv_654: n_907  <= TRANSPORT NOT a_LC3_D22  ;
inv_655: n_908  <= TRANSPORT NOT a_N2353  ;
delay_656: n_909  <= TRANSPORT dbin(6)  ;
and2_657: n_910 <=  n_911  AND n_912;
delay_658: n_911  <= TRANSPORT a_N2353  ;
delay_659: n_912  <= TRANSPORT a_SCH0BWORDOUT_F14_G  ;
and2_660: n_913 <=  n_914  AND n_915;
delay_661: n_914  <= TRANSPORT a_LC3_D22  ;
delay_662: n_915  <= TRANSPORT a_SCH0BWORDOUT_F14_G  ;
and1_663: n_916 <=  gnd;
delay_664: n_917  <= TRANSPORT clk  ;
filter_665: FILTER_a8237

    PORT MAP (IN1 => n_917, Y => a_SCH0BWORDOUT_F14_G_aCLK);
delay_666: a_LC1_C22  <= TRANSPORT a_EQ024  ;
xor2_667: a_EQ024 <=  n_921  XOR n_935;
or3_668: n_921 <=  n_922  OR n_927  OR n_931;
and2_669: n_922 <=  n_923  AND n_925;
inv_670: n_923  <= TRANSPORT NOT a_N3554  ;
delay_671: n_925  <= TRANSPORT a_N3556  ;
and2_672: n_927 <=  n_928  AND n_929;
inv_673: n_928  <= TRANSPORT NOT a_N3554  ;
delay_674: n_929  <= TRANSPORT a_N3555  ;
and3_675: n_931 <=  n_932  AND n_933  AND n_934;
delay_676: n_932  <= TRANSPORT a_N3554  ;
inv_677: n_933  <= TRANSPORT NOT a_N3555  ;
inv_678: n_934  <= TRANSPORT NOT a_N3556  ;
and1_679: n_935 <=  gnd;
delay_680: a_LC4_A3  <= TRANSPORT a_EQ192  ;
xor2_681: a_EQ192 <=  n_938  XOR n_945;
or3_682: n_938 <=  n_939  OR n_941  OR n_943;
and1_683: n_939 <=  n_940;
inv_684: n_940  <= TRANSPORT NOT ain(3)  ;
and1_685: n_941 <=  n_942;
inv_686: n_942  <= TRANSPORT NOT ain(2)  ;
and1_687: n_943 <=  n_944;
delay_688: n_944  <= TRANSPORT ain(1)  ;
and1_689: n_945 <=  gnd;
delay_690: a_N2563_aNOT  <= TRANSPORT a_EQ616  ;
xor2_691: a_EQ616 <=  n_948  XOR n_955;
or3_692: n_948 <=  n_949  OR n_951  OR n_953;
and1_693: n_949 <=  n_950;
inv_694: n_950  <= TRANSPORT NOT ain(0)  ;
and1_695: n_951 <=  n_952;
delay_696: n_952  <= TRANSPORT a_LC4_A3  ;
and1_697: n_953 <=  n_954;
delay_698: n_954  <= TRANSPORT a_N87  ;
and1_699: n_955 <=  gnd;
delay_700: a_N70  <= TRANSPORT a_N70_aIN  ;
xor2_701: a_N70_aIN <=  n_958  XOR n_968;
or1_702: n_958 <=  n_959;
and4_703: n_959 <=  n_960  AND n_962  AND n_964  AND n_966;
delay_704: n_960  <= TRANSPORT a_N820  ;
delay_705: n_962  <= TRANSPORT a_N822  ;
inv_706: n_964  <= TRANSPORT NOT a_N821  ;
inv_707: n_966  <= TRANSPORT NOT a_N823  ;
and1_708: n_968 <=  gnd;
delay_709: a_N71_aNOT  <= TRANSPORT a_EQ190  ;
xor2_710: a_EQ190 <=  n_971  XOR n_980;
or4_711: n_971 <=  n_972  OR n_974  OR n_976  OR n_978;
and1_712: n_972 <=  n_973;
inv_713: n_973  <= TRANSPORT NOT a_N820  ;
and1_714: n_974 <=  n_975;
inv_715: n_975  <= TRANSPORT NOT a_N821  ;
and1_716: n_976 <=  n_977;
delay_717: n_977  <= TRANSPORT a_N823  ;
and1_718: n_978 <=  n_979;
inv_719: n_979  <= TRANSPORT NOT a_N822  ;
and1_720: n_980 <=  gnd;
delay_721: a_LC1_B23_aNOT  <= TRANSPORT a_EQ574  ;
xor2_722: a_EQ574 <=  n_983  XOR n_990;
or3_723: n_983 <=  n_984  OR n_986  OR n_988;
and1_724: n_984 <=  n_985;
inv_725: n_985  <= TRANSPORT NOT a_N821  ;
and1_726: n_986 <=  n_987;
delay_727: n_987  <= TRANSPORT a_N823  ;
and1_728: n_988 <=  n_989;
inv_729: n_989  <= TRANSPORT NOT a_N822  ;
and1_730: n_990 <=  gnd;
delay_731: a_N2361  <= TRANSPORT a_EQ562  ;
xor2_732: a_EQ562 <=  n_993  XOR n_998;
or2_733: n_993 <=  n_994  OR n_996;
and1_734: n_994 <=  n_995;
delay_735: n_995  <= TRANSPORT a_N820  ;
and1_736: n_996 <=  n_997;
delay_737: n_997  <= TRANSPORT a_LC1_B23_aNOT  ;
and1_738: n_998 <=  gnd;
delay_739: a_N1584  <= TRANSPORT a_EQ472  ;
xor2_740: a_EQ472 <=  n_1001  XOR n_1008;
or3_741: n_1001 <=  n_1002  OR n_1004  OR n_1006;
and1_742: n_1002 <=  n_1003;
delay_743: n_1003  <= TRANSPORT a_N70  ;
and1_744: n_1004 <=  n_1005;
inv_745: n_1005  <= TRANSPORT NOT a_N71_aNOT  ;
and1_746: n_1006 <=  n_1007;
inv_747: n_1007  <= TRANSPORT NOT a_N2361  ;
and1_748: n_1008 <=  gnd;
delay_749: a_N2557  <= TRANSPORT a_N2557_aIN  ;
xor2_750: a_N2557_aIN <=  n_1011  XOR n_1015;
or1_751: n_1011 <=  n_1012;
and2_752: n_1012 <=  n_1013  AND n_1014;
delay_753: n_1013  <= TRANSPORT a_N2563_aNOT  ;
delay_754: n_1014  <= TRANSPORT a_N1584  ;
and1_755: n_1015 <=  gnd;
delay_756: a_N1164_aNOT  <= TRANSPORT a_EQ374  ;
xor2_757: a_EQ374 <=  n_1018  XOR n_1025;
or2_758: n_1018 <=  n_1019  OR n_1022;
and2_759: n_1019 <=  n_1020  AND n_1021;
inv_760: n_1020  <= TRANSPORT NOT a_LC1_C22  ;
delay_761: n_1021  <= TRANSPORT a_N2557  ;
and2_762: n_1022 <=  n_1023  AND n_1024;
inv_763: n_1023  <= TRANSPORT NOT a_N2557  ;
delay_764: n_1024  <= TRANSPORT a_N3554  ;
and1_765: n_1025 <=  gnd;
delay_766: a_N2598_aNOT  <= TRANSPORT a_EQ647  ;
xor2_767: a_EQ647 <=  n_1028  XOR n_1035;
or2_768: n_1028 <=  n_1029  OR n_1032;
and1_769: n_1029 <=  n_1030;
delay_770: n_1030  <= TRANSPORT a_SCHANNEL_F1_G  ;
and1_771: n_1032 <=  n_1033;
delay_772: n_1033  <= TRANSPORT a_SCHANNEL_F0_G  ;
and1_773: n_1035 <=  gnd;
delay_774: a_N2591  <= TRANSPORT a_N2591_aIN  ;
xor2_775: a_N2591_aIN <=  n_1038  XOR n_1043;
or1_776: n_1038 <=  n_1039;
and2_777: n_1039 <=  n_1040  AND n_1041;
inv_778: n_1040  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_779: n_1041  <= TRANSPORT a_SCOMMANDREG_F0_G  ;
and1_780: n_1043 <=  gnd;
delay_781: a_N2531  <= TRANSPORT a_N2531_aIN  ;
xor2_782: a_N2531_aIN <=  n_1046  XOR n_1050;
or1_783: n_1046 <=  n_1047;
and2_784: n_1047 <=  n_1048  AND n_1049;
delay_785: n_1048  <= TRANSPORT a_N2557  ;
delay_786: n_1049  <= TRANSPORT a_N2591  ;
and1_787: n_1050 <=  gnd;
delay_788: a_N2374  <= TRANSPORT a_EQ568  ;
xor2_789: a_EQ568 <=  n_1053  XOR n_1062;
or4_790: n_1053 <=  n_1054  OR n_1056  OR n_1058  OR n_1060;
and1_791: n_1054 <=  n_1055;
inv_792: n_1055  <= TRANSPORT NOT a_N820  ;
and1_793: n_1056 <=  n_1057;
inv_794: n_1057  <= TRANSPORT NOT a_N823  ;
and1_795: n_1058 <=  n_1059;
inv_796: n_1059  <= TRANSPORT NOT a_N822  ;
and1_797: n_1060 <=  n_1061;
delay_798: n_1061  <= TRANSPORT a_N821  ;
and1_799: n_1062 <=  gnd;
delay_800: a_N2408_aNOT  <= TRANSPORT a_EQ579  ;
xor2_801: a_EQ579 <=  n_1065  XOR n_1078;
or4_802: n_1065 <=  n_1066  OR n_1069  OR n_1072  OR n_1075;
and2_803: n_1066 <=  n_1067  AND n_1068;
delay_804: n_1067  <= TRANSPORT a_N822  ;
inv_805: n_1068  <= TRANSPORT NOT a_N821  ;
and2_806: n_1069 <=  n_1070  AND n_1071;
inv_807: n_1070  <= TRANSPORT NOT a_N822  ;
delay_808: n_1071  <= TRANSPORT a_N823  ;
and2_809: n_1072 <=  n_1073  AND n_1074;
inv_810: n_1073  <= TRANSPORT NOT a_N820  ;
inv_811: n_1074  <= TRANSPORT NOT a_N823  ;
and2_812: n_1075 <=  n_1076  AND n_1077;
delay_813: n_1076  <= TRANSPORT a_N821  ;
inv_814: n_1077  <= TRANSPORT NOT a_N823  ;
and1_815: n_1078 <=  gnd;
delay_816: a_N68_aNOT  <= TRANSPORT a_EQ188  ;
xor2_817: a_EQ188 <=  n_1081  XOR n_1090;
or4_818: n_1081 <=  n_1082  OR n_1084  OR n_1086  OR n_1088;
and1_819: n_1082 <=  n_1083;
delay_820: n_1083  <= TRANSPORT a_N820  ;
and1_821: n_1084 <=  n_1085;
inv_822: n_1085  <= TRANSPORT NOT a_N823  ;
and1_823: n_1086 <=  n_1087;
inv_824: n_1087  <= TRANSPORT NOT a_N822  ;
and1_825: n_1088 <=  n_1089;
delay_826: n_1089  <= TRANSPORT a_N821  ;
and1_827: n_1090 <=  gnd;
delay_828: a_LC4_B25_aNOT  <= TRANSPORT a_LC4_B25_aNOT_aIN  ;
xor2_829: a_LC4_B25_aNOT_aIN <=  n_1093  XOR n_1097;
or1_830: n_1093 <=  n_1094;
and2_831: n_1094 <=  n_1095  AND n_1096;
delay_832: n_1095  <= TRANSPORT a_N2408_aNOT  ;
delay_833: n_1096  <= TRANSPORT a_N68_aNOT  ;
and1_834: n_1097 <=  gnd;
delay_835: a_N67_aNOT  <= TRANSPORT a_EQ187  ;
xor2_836: a_EQ187 <=  n_1100  XOR n_1109;
or4_837: n_1100 <=  n_1101  OR n_1103  OR n_1105  OR n_1107;
and1_838: n_1101 <=  n_1102;
inv_839: n_1102  <= TRANSPORT NOT a_N823  ;
and1_840: n_1103 <=  n_1104;
delay_841: n_1104  <= TRANSPORT a_N820  ;
and1_842: n_1105 <=  n_1106;
delay_843: n_1106  <= TRANSPORT a_N822  ;
and1_844: n_1107 <=  n_1108;
inv_845: n_1108  <= TRANSPORT NOT a_N821  ;
and1_846: n_1109 <=  gnd;
delay_847: a_N2356  <= TRANSPORT a_EQ559  ;
xor2_848: a_EQ559 <=  n_1112  XOR n_1121;
or4_849: n_1112 <=  n_1113  OR n_1115  OR n_1117  OR n_1119;
and1_850: n_1113 <=  n_1114;
delay_851: n_1114  <= TRANSPORT a_N823  ;
and1_852: n_1115 <=  n_1116;
delay_853: n_1116  <= TRANSPORT a_N820  ;
and1_854: n_1117 <=  n_1118;
delay_855: n_1118  <= TRANSPORT a_N822  ;
and1_856: n_1119 <=  n_1120;
inv_857: n_1120  <= TRANSPORT NOT a_N821  ;
and1_858: n_1121 <=  gnd;
delay_859: a_N1592  <= TRANSPORT a_N1592_aIN  ;
xor2_860: a_N1592_aIN <=  n_1124  XOR n_1129;
or1_861: n_1124 <=  n_1125;
and3_862: n_1125 <=  n_1126  AND n_1127  AND n_1128;
delay_863: n_1126  <= TRANSPORT a_N2361  ;
delay_864: n_1127  <= TRANSPORT a_N67_aNOT  ;
delay_865: n_1128  <= TRANSPORT a_N2356  ;
and1_866: n_1129 <=  gnd;
delay_867: a_N1566  <= TRANSPORT a_EQ465  ;
xor2_868: a_EQ465 <=  n_1132  XOR n_1139;
or3_869: n_1132 <=  n_1133  OR n_1135  OR n_1137;
and1_870: n_1133 <=  n_1134;
delay_871: n_1134  <= TRANSPORT a_N820  ;
and1_872: n_1135 <=  n_1136;
delay_873: n_1136  <= TRANSPORT a_N822  ;
and1_874: n_1137 <=  n_1138;
delay_875: n_1138  <= TRANSPORT a_N821  ;
and1_876: n_1139 <=  gnd;
delay_877: a_N2358  <= TRANSPORT a_EQ560  ;
xor2_878: a_EQ560 <=  n_1142  XOR n_1151;
or4_879: n_1142 <=  n_1143  OR n_1145  OR n_1147  OR n_1149;
and1_880: n_1143 <=  n_1144;
delay_881: n_1144  <= TRANSPORT a_N820  ;
and1_882: n_1145 <=  n_1146;
delay_883: n_1146  <= TRANSPORT a_N823  ;
and1_884: n_1147 <=  n_1148;
inv_885: n_1148  <= TRANSPORT NOT a_N822  ;
and1_886: n_1149 <=  n_1150;
delay_887: n_1150  <= TRANSPORT a_N821  ;
and1_888: n_1151 <=  gnd;
delay_889: a_LC8_B20  <= TRANSPORT a_EQ476  ;
xor2_890: a_EQ476 <=  n_1154  XOR n_1164;
or3_891: n_1154 <=  n_1155  OR n_1158  OR n_1161;
and2_892: n_1155 <=  n_1156  AND n_1157;
delay_893: n_1156  <= TRANSPORT a_N2563_aNOT  ;
inv_894: n_1157  <= TRANSPORT NOT a_N820  ;
and2_895: n_1158 <=  n_1159  AND n_1160;
delay_896: n_1159  <= TRANSPORT a_N2563_aNOT  ;
delay_897: n_1160  <= TRANSPORT a_N822  ;
and2_898: n_1161 <=  n_1162  AND n_1163;
delay_899: n_1162  <= TRANSPORT a_N2563_aNOT  ;
inv_900: n_1163  <= TRANSPORT NOT a_N821  ;
and1_901: n_1164 <=  gnd;
delay_902: a_N1588  <= TRANSPORT a_N1588_aIN  ;
xor2_903: a_N1588_aIN <=  n_1167  XOR n_1172;
or1_904: n_1167 <=  n_1168;
and3_905: n_1168 <=  n_1169  AND n_1170  AND n_1171;
delay_906: n_1169  <= TRANSPORT a_N1566  ;
delay_907: n_1170  <= TRANSPORT a_N2358  ;
delay_908: n_1171  <= TRANSPORT a_LC8_B20  ;
and1_909: n_1172 <=  gnd;
delay_910: a_N88_aNOT  <= TRANSPORT a_EQ197  ;
xor2_911: a_EQ197 <=  n_1175  XOR n_1180;
or2_912: n_1175 <=  n_1176  OR n_1178;
and1_913: n_1176 <=  n_1177;
delay_914: n_1177  <= TRANSPORT a_SCHANNEL_F1_G  ;
and1_915: n_1178 <=  n_1179;
inv_916: n_1179  <= TRANSPORT NOT a_SCHANNEL_F0_G  ;
and1_917: n_1180 <=  gnd;
delay_918: a_N2377  <= TRANSPORT a_EQ570  ;
xor2_919: a_EQ570 <=  n_1183  XOR n_1188;
or2_920: n_1183 <=  n_1184  OR n_1186;
and1_921: n_1184 <=  n_1185;
inv_922: n_1185  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and1_923: n_1186 <=  n_1187;
inv_924: n_1187  <= TRANSPORT NOT a_SCHANNEL_F0_G  ;
and1_925: n_1188 <=  gnd;
delay_926: a_LC4_E22  <= TRANSPORT a_EQ580  ;
xor2_927: a_EQ580 <=  n_1191  XOR n_1200;
or2_928: n_1191 <=  n_1192  OR n_1196;
and2_929: n_1192 <=  n_1193  AND n_1194;
inv_930: n_1193  <= TRANSPORT NOT a_N88_aNOT  ;
delay_931: n_1194  <= TRANSPORT a_SCH1MODEREG_F1_G  ;
and2_932: n_1196 <=  n_1197  AND n_1198;
inv_933: n_1197  <= TRANSPORT NOT a_N2377  ;
delay_934: n_1198  <= TRANSPORT a_SCH3MODEREG_F1_G  ;
and1_935: n_1200 <=  gnd;
delay_936: a_N2376  <= TRANSPORT a_EQ569  ;
xor2_937: a_EQ569 <=  n_1203  XOR n_1208;
or2_938: n_1203 <=  n_1204  OR n_1206;
and1_939: n_1204 <=  n_1205;
inv_940: n_1205  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and1_941: n_1206 <=  n_1207;
delay_942: n_1207  <= TRANSPORT a_SCHANNEL_F0_G  ;
and1_943: n_1208 <=  gnd;
delay_944: a_LC6_E22  <= TRANSPORT a_EQ582  ;
xor2_945: a_EQ582 <=  n_1211  XOR n_1226;
or4_946: n_1211 <=  n_1212  OR n_1217  OR n_1220  OR n_1223;
and2_947: n_1212 <=  n_1213  AND n_1215;
inv_948: n_1213  <= TRANSPORT NOT a_SCH2MODEREG_F0_G  ;
inv_949: n_1215  <= TRANSPORT NOT a_SCH1MODEREG_F0_G  ;
and2_950: n_1217 <=  n_1218  AND n_1219;
delay_951: n_1218  <= TRANSPORT a_N88_aNOT  ;
inv_952: n_1219  <= TRANSPORT NOT a_SCH2MODEREG_F0_G  ;
and2_953: n_1220 <=  n_1221  AND n_1222;
delay_954: n_1221  <= TRANSPORT a_N2376  ;
inv_955: n_1222  <= TRANSPORT NOT a_SCH1MODEREG_F0_G  ;
and2_956: n_1223 <=  n_1224  AND n_1225;
delay_957: n_1224  <= TRANSPORT a_N88_aNOT  ;
delay_958: n_1225  <= TRANSPORT a_N2376  ;
and1_959: n_1226 <=  gnd;
delay_960: a_LC5_E22  <= TRANSPORT a_EQ583  ;
xor2_961: a_EQ583 <=  n_1229  XOR n_1244;
or4_962: n_1229 <=  n_1230  OR n_1235  OR n_1238  OR n_1241;
and2_963: n_1230 <=  n_1231  AND n_1233;
inv_964: n_1231  <= TRANSPORT NOT a_SCH0MODEREG_F0_G  ;
inv_965: n_1233  <= TRANSPORT NOT a_SCH3MODEREG_F0_G  ;
and2_966: n_1235 <=  n_1236  AND n_1237;
delay_967: n_1236  <= TRANSPORT a_N2377  ;
inv_968: n_1237  <= TRANSPORT NOT a_SCH0MODEREG_F0_G  ;
and2_969: n_1238 <=  n_1239  AND n_1240;
delay_970: n_1239  <= TRANSPORT a_N2598_aNOT  ;
inv_971: n_1240  <= TRANSPORT NOT a_SCH3MODEREG_F0_G  ;
and2_972: n_1241 <=  n_1242  AND n_1243;
delay_973: n_1242  <= TRANSPORT a_N2598_aNOT  ;
delay_974: n_1243  <= TRANSPORT a_N2377  ;
and1_975: n_1244 <=  gnd;
delay_976: a_LC6_E10  <= TRANSPORT a_EQ581  ;
xor2_977: a_EQ581 <=  n_1247  XOR n_1256;
or2_978: n_1247 <=  n_1248  OR n_1252;
and2_979: n_1248 <=  n_1249  AND n_1250;
inv_980: n_1249  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_981: n_1250  <= TRANSPORT a_SCH0MODEREG_F1_G  ;
and2_982: n_1252 <=  n_1253  AND n_1254;
inv_983: n_1253  <= TRANSPORT NOT a_N2376  ;
delay_984: n_1254  <= TRANSPORT a_SCH2MODEREG_F1_G  ;
and1_985: n_1256 <=  gnd;
delay_986: a_N1589  <= TRANSPORT a_EQ478  ;
xor2_987: a_EQ478 <=  n_1259  XOR n_1268;
or2_988: n_1259 <=  n_1260  OR n_1264;
and3_989: n_1260 <=  n_1261  AND n_1262  AND n_1263;
delay_990: n_1261  <= TRANSPORT a_LC4_E22  ;
delay_991: n_1262  <= TRANSPORT a_LC6_E22  ;
delay_992: n_1263  <= TRANSPORT a_LC5_E22  ;
and3_993: n_1264 <=  n_1265  AND n_1266  AND n_1267;
delay_994: n_1265  <= TRANSPORT a_LC6_E22  ;
delay_995: n_1266  <= TRANSPORT a_LC5_E22  ;
delay_996: n_1267  <= TRANSPORT a_LC6_E10  ;
and1_997: n_1268 <=  gnd;
delay_998: a_N1580_aNOT  <= TRANSPORT a_EQ468  ;
xor2_999: a_EQ468 <=  n_1271  XOR n_1280;
or2_1000: n_1271 <=  n_1272  OR n_1276;
and3_1001: n_1272 <=  n_1273  AND n_1274  AND n_1275;
delay_1002: n_1273  <= TRANSPORT a_N71_aNOT  ;
delay_1003: n_1274  <= TRANSPORT a_N1592  ;
delay_1004: n_1275  <= TRANSPORT a_N1588  ;
and3_1005: n_1276 <=  n_1277  AND n_1278  AND n_1279;
delay_1006: n_1277  <= TRANSPORT a_N71_aNOT  ;
delay_1007: n_1278  <= TRANSPORT a_N1588  ;
delay_1008: n_1279  <= TRANSPORT a_N1589  ;
and1_1009: n_1280 <=  gnd;
delay_1010: a_SNMEMR_aNOT  <= TRANSPORT a_SNMEMR_aNOT_aIN  ;
xor2_1011: a_SNMEMR_aNOT_aIN <=  n_1282  XOR n_1287;
or1_1012: n_1282 <=  n_1283;
and3_1013: n_1283 <=  n_1284  AND n_1285  AND n_1286;
delay_1014: n_1284  <= TRANSPORT a_N2374  ;
delay_1015: n_1285  <= TRANSPORT a_LC4_B25_aNOT  ;
delay_1016: n_1286  <= TRANSPORT a_N1580_aNOT  ;
and1_1017: n_1287 <=  gnd;
delay_1018: a_N1180  <= TRANSPORT a_EQ385  ;
xor2_1019: a_EQ385 <=  n_1290  XOR n_1299;
or2_1020: n_1290 <=  n_1291  OR n_1295;
and2_1021: n_1291 <=  n_1292  AND n_1293;
delay_1022: n_1292  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_1023: n_1293  <= TRANSPORT a_SCH1WRDCNTREG_F2_G  ;
and2_1024: n_1295 <=  n_1296  AND n_1297;
inv_1025: n_1296  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_1026: n_1297  <= TRANSPORT a_SCH0WRDCNTREG_F2_G  ;
and1_1027: n_1299 <=  gnd;
delay_1028: a_LC4_C6  <= TRANSPORT a_EQ386  ;
xor2_1029: a_EQ386 <=  n_1302  XOR n_1309;
or2_1030: n_1302 <=  n_1303  OR n_1306;
and2_1031: n_1303 <=  n_1304  AND n_1305;
delay_1032: n_1304  <= TRANSPORT a_N1164_aNOT  ;
inv_1033: n_1305  <= TRANSPORT NOT a_N2531  ;
and2_1034: n_1306 <=  n_1307  AND n_1308;
delay_1035: n_1307  <= TRANSPORT a_N2531  ;
delay_1036: n_1308  <= TRANSPORT a_N1180  ;
and1_1037: n_1309 <=  gnd;
delay_1038: a_LC2_C6  <= TRANSPORT a_EQ384  ;
xor2_1039: a_EQ384 <=  n_1312  XOR n_1321;
or2_1040: n_1312 <=  n_1313  OR n_1317;
and2_1041: n_1313 <=  n_1314  AND n_1315;
inv_1042: n_1314  <= TRANSPORT NOT a_N2376  ;
delay_1043: n_1315  <= TRANSPORT a_SCH2WRDCNTREG_F2_G  ;
and2_1044: n_1317 <=  n_1318  AND n_1319;
inv_1045: n_1318  <= TRANSPORT NOT a_N2377  ;
delay_1046: n_1319  <= TRANSPORT a_SCH3WRDCNTREG_F2_G  ;
and1_1047: n_1321 <=  gnd;
delay_1048: a_LC1_C6  <= TRANSPORT a_EQ383  ;
xor2_1049: a_EQ383 <=  n_1324  XOR n_1331;
or2_1050: n_1324 <=  n_1325  OR n_1328;
and2_1051: n_1325 <=  n_1326  AND n_1327;
inv_1052: n_1326  <= TRANSPORT NOT a_N88_aNOT  ;
delay_1053: n_1327  <= TRANSPORT a_SCH1WRDCNTREG_F2_G  ;
and2_1054: n_1328 <=  n_1329  AND n_1330;
inv_1055: n_1329  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_1056: n_1330  <= TRANSPORT a_SCH0WRDCNTREG_F2_G  ;
and1_1057: n_1331 <=  gnd;
dff_1058: DFF_a8237

    PORT MAP ( D => a_EQ850, CLK => a_N3554_aCLK, CLRN => a_N3554_aCLRN, PRN => vcc,
          Q => a_N3554);
inv_1059: a_N3554_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1060: a_EQ850 <=  n_1338  XOR n_1349;
or3_1061: n_1338 <=  n_1339  OR n_1343  OR n_1346;
and2_1062: n_1339 <=  n_1340  AND n_1341;
delay_1063: n_1340  <= TRANSPORT a_LC4_C6  ;
inv_1064: n_1341  <= TRANSPORT NOT startdma  ;
and2_1065: n_1343 <=  n_1344  AND n_1345;
delay_1066: n_1344  <= TRANSPORT a_LC2_C6  ;
delay_1067: n_1345  <= TRANSPORT startdma  ;
and2_1068: n_1346 <=  n_1347  AND n_1348;
delay_1069: n_1347  <= TRANSPORT a_LC1_C6  ;
delay_1070: n_1348  <= TRANSPORT startdma  ;
and1_1071: n_1349 <=  gnd;
delay_1072: n_1350  <= TRANSPORT clk  ;
filter_1073: FILTER_a8237

    PORT MAP (IN1 => n_1350, Y => a_N3554_aCLK);
delay_1074: a_LC7_C22  <= TRANSPORT a_EQ023  ;
xor2_1075: a_EQ023 <=  n_1354  XOR n_1361;
or2_1076: n_1354 <=  n_1355  OR n_1358;
and2_1077: n_1355 <=  n_1356  AND n_1357;
inv_1078: n_1356  <= TRANSPORT NOT a_N3555  ;
delay_1079: n_1357  <= TRANSPORT a_N3556  ;
and2_1080: n_1358 <=  n_1359  AND n_1360;
delay_1081: n_1359  <= TRANSPORT a_N3555  ;
inv_1082: n_1360  <= TRANSPORT NOT a_N3556  ;
and1_1083: n_1361 <=  gnd;
delay_1084: a_LC4_C27  <= TRANSPORT a_EQ361  ;
xor2_1085: a_EQ361 <=  n_1364  XOR n_1372;
or2_1086: n_1364 <=  n_1365  OR n_1369;
and3_1087: n_1365 <=  n_1366  AND n_1367  AND n_1368;
delay_1088: n_1366  <= TRANSPORT a_N2557  ;
inv_1089: n_1367  <= TRANSPORT NOT a_N2531  ;
inv_1090: n_1368  <= TRANSPORT NOT a_LC7_C22  ;
and2_1091: n_1369 <=  n_1370  AND n_1371;
inv_1092: n_1370  <= TRANSPORT NOT a_N2557  ;
delay_1093: n_1371  <= TRANSPORT a_N3555  ;
and1_1094: n_1372 <=  gnd;
delay_1095: a_LC6_C27  <= TRANSPORT a_EQ363  ;
xor2_1096: a_EQ363 <=  n_1375  XOR n_1384;
or2_1097: n_1375 <=  n_1376  OR n_1380;
and2_1098: n_1376 <=  n_1377  AND n_1378;
inv_1099: n_1377  <= TRANSPORT NOT a_N88_aNOT  ;
delay_1100: n_1378  <= TRANSPORT a_SCH1WRDCNTREG_F1_G  ;
and2_1101: n_1380 <=  n_1381  AND n_1382;
inv_1102: n_1381  <= TRANSPORT NOT a_N2377  ;
delay_1103: n_1382  <= TRANSPORT a_SCH3WRDCNTREG_F1_G  ;
and1_1104: n_1384 <=  gnd;
delay_1105: a_LC2_C27  <= TRANSPORT a_EQ364  ;
xor2_1106: a_EQ364 <=  n_1387  XOR n_1396;
or2_1107: n_1387 <=  n_1388  OR n_1392;
and2_1108: n_1388 <=  n_1389  AND n_1390;
inv_1109: n_1389  <= TRANSPORT NOT a_N2376  ;
delay_1110: n_1390  <= TRANSPORT a_SCH2WRDCNTREG_F1_G  ;
and2_1111: n_1392 <=  n_1393  AND n_1394;
inv_1112: n_1393  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_1113: n_1394  <= TRANSPORT a_SCH0WRDCNTREG_F1_G  ;
and1_1114: n_1396 <=  gnd;
delay_1115: a_N1139  <= TRANSPORT a_EQ365  ;
xor2_1116: a_EQ365 <=  n_1399  XOR n_1406;
or3_1117: n_1399 <=  n_1400  OR n_1402  OR n_1404;
and1_1118: n_1400 <=  n_1401;
delay_1119: n_1401  <= TRANSPORT a_LC6_C27  ;
and1_1120: n_1402 <=  n_1403;
inv_1121: n_1403  <= TRANSPORT NOT startdma  ;
and1_1122: n_1404 <=  n_1405;
delay_1123: n_1405  <= TRANSPORT a_LC2_C27  ;
and1_1124: n_1406 <=  gnd;
delay_1125: a_LC5_C27  <= TRANSPORT a_EQ362  ;
xor2_1126: a_EQ362 <=  n_1409  XOR n_1418;
or2_1127: n_1409 <=  n_1410  OR n_1414;
and3_1128: n_1410 <=  n_1411  AND n_1412  AND n_1413;
delay_1129: n_1411  <= TRANSPORT a_N2531  ;
delay_1130: n_1412  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_1131: n_1413  <= TRANSPORT a_SCH1WRDCNTREG_F1_G  ;
and3_1132: n_1414 <=  n_1415  AND n_1416  AND n_1417;
delay_1133: n_1415  <= TRANSPORT a_N2531  ;
inv_1134: n_1416  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_1135: n_1417  <= TRANSPORT a_SCH0WRDCNTREG_F1_G  ;
and1_1136: n_1418 <=  gnd;
dff_1137: DFF_a8237

    PORT MAP ( D => a_EQ851, CLK => a_N3555_aCLK, CLRN => a_N3555_aCLRN, PRN => vcc,
          Q => a_N3555);
inv_1138: a_N3555_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1139: a_EQ851 <=  n_1425  XOR n_1435;
or3_1140: n_1425 <=  n_1426  OR n_1429  OR n_1432;
and2_1141: n_1426 <=  n_1427  AND n_1428;
delay_1142: n_1427  <= TRANSPORT a_LC4_C27  ;
delay_1143: n_1428  <= TRANSPORT a_N1139  ;
and2_1144: n_1429 <=  n_1430  AND n_1431;
delay_1145: n_1430  <= TRANSPORT a_N1139  ;
delay_1146: n_1431  <= TRANSPORT startdma  ;
and2_1147: n_1432 <=  n_1433  AND n_1434;
delay_1148: n_1433  <= TRANSPORT a_N1139  ;
delay_1149: n_1434  <= TRANSPORT a_LC5_C27  ;
and1_1150: n_1435 <=  gnd;
delay_1151: n_1436  <= TRANSPORT clk  ;
filter_1152: FILTER_a8237

    PORT MAP (IN1 => n_1436, Y => a_N3555_aCLK);
delay_1153: a_LC1_C21  <= TRANSPORT a_EQ025  ;
xor2_1154: a_EQ025 <=  n_1440  XOR n_1456;
or4_1155: n_1440 <=  n_1441  OR n_1445  OR n_1448  OR n_1451;
and2_1156: n_1441 <=  n_1442  AND n_1443;
delay_1157: n_1442  <= TRANSPORT a_N3554  ;
inv_1158: n_1443  <= TRANSPORT NOT a_N3553  ;
and2_1159: n_1445 <=  n_1446  AND n_1447;
inv_1160: n_1446  <= TRANSPORT NOT a_N3553  ;
delay_1161: n_1447  <= TRANSPORT a_N3556  ;
and2_1162: n_1448 <=  n_1449  AND n_1450;
delay_1163: n_1449  <= TRANSPORT a_N3555  ;
inv_1164: n_1450  <= TRANSPORT NOT a_N3553  ;
and4_1165: n_1451 <=  n_1452  AND n_1453  AND n_1454  AND n_1455;
inv_1166: n_1452  <= TRANSPORT NOT a_N3554  ;
inv_1167: n_1453  <= TRANSPORT NOT a_N3555  ;
delay_1168: n_1454  <= TRANSPORT a_N3553  ;
inv_1169: n_1455  <= TRANSPORT NOT a_N3556  ;
and1_1170: n_1456 <=  gnd;
delay_1171: a_LC7_C15  <= TRANSPORT a_EQ253  ;
xor2_1172: a_EQ253 <=  n_1459  XOR n_1466;
or2_1173: n_1459 <=  n_1460  OR n_1463;
and2_1174: n_1460 <=  n_1461  AND n_1462;
inv_1175: n_1461  <= TRANSPORT NOT a_N2557  ;
delay_1176: n_1462  <= TRANSPORT a_N3553  ;
and2_1177: n_1463 <=  n_1464  AND n_1465;
delay_1178: n_1464  <= TRANSPORT a_N2557  ;
inv_1179: n_1465  <= TRANSPORT NOT a_LC1_C21  ;
and1_1180: n_1466 <=  gnd;
delay_1181: a_LC5_C15  <= TRANSPORT a_EQ254  ;
xor2_1182: a_EQ254 <=  n_1469  XOR n_1478;
or2_1183: n_1469 <=  n_1470  OR n_1474;
and2_1184: n_1470 <=  n_1471  AND n_1472;
delay_1185: n_1471  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_1186: n_1472  <= TRANSPORT a_SCH1WRDCNTREG_F3_G  ;
and2_1187: n_1474 <=  n_1475  AND n_1476;
inv_1188: n_1475  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_1189: n_1476  <= TRANSPORT a_SCH0WRDCNTREG_F3_G  ;
and1_1190: n_1478 <=  gnd;
delay_1191: a_N491_aNOT  <= TRANSPORT a_EQ255  ;
xor2_1192: a_EQ255 <=  n_1481  XOR n_1488;
or2_1193: n_1481 <=  n_1482  OR n_1485;
and2_1194: n_1482 <=  n_1483  AND n_1484;
inv_1195: n_1483  <= TRANSPORT NOT a_N2531  ;
delay_1196: n_1484  <= TRANSPORT a_LC7_C15  ;
and2_1197: n_1485 <=  n_1486  AND n_1487;
delay_1198: n_1486  <= TRANSPORT a_N2531  ;
delay_1199: n_1487  <= TRANSPORT a_LC5_C15  ;
and1_1200: n_1488 <=  gnd;
delay_1201: a_LC5_C14  <= TRANSPORT a_EQ257  ;
xor2_1202: a_EQ257 <=  n_1491  XOR n_1500;
or2_1203: n_1491 <=  n_1492  OR n_1496;
and2_1204: n_1492 <=  n_1493  AND n_1494;
inv_1205: n_1493  <= TRANSPORT NOT a_N2377  ;
delay_1206: n_1494  <= TRANSPORT a_SCH3WRDCNTREG_F3_G  ;
and2_1207: n_1496 <=  n_1497  AND n_1498;
inv_1208: n_1497  <= TRANSPORT NOT a_N2376  ;
delay_1209: n_1498  <= TRANSPORT a_SCH2WRDCNTREG_F3_G  ;
and1_1210: n_1500 <=  gnd;
delay_1211: a_LC1_C15  <= TRANSPORT a_EQ256  ;
xor2_1212: a_EQ256 <=  n_1503  XOR n_1510;
or2_1213: n_1503 <=  n_1504  OR n_1507;
and2_1214: n_1504 <=  n_1505  AND n_1506;
inv_1215: n_1505  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_1216: n_1506  <= TRANSPORT a_SCH0WRDCNTREG_F3_G  ;
and2_1217: n_1507 <=  n_1508  AND n_1509;
inv_1218: n_1508  <= TRANSPORT NOT a_N88_aNOT  ;
delay_1219: n_1509  <= TRANSPORT a_SCH1WRDCNTREG_F3_G  ;
and1_1220: n_1510 <=  gnd;
dff_1221: DFF_a8237

    PORT MAP ( D => a_EQ849, CLK => a_N3553_aCLK, CLRN => a_N3553_aCLRN, PRN => vcc,
          Q => a_N3553);
inv_1222: a_N3553_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1223: a_EQ849 <=  n_1517  XOR n_1527;
or3_1224: n_1517 <=  n_1518  OR n_1521  OR n_1524;
and2_1225: n_1518 <=  n_1519  AND n_1520;
delay_1226: n_1519  <= TRANSPORT a_N491_aNOT  ;
inv_1227: n_1520  <= TRANSPORT NOT startdma  ;
and2_1228: n_1521 <=  n_1522  AND n_1523;
delay_1229: n_1522  <= TRANSPORT a_LC5_C14  ;
delay_1230: n_1523  <= TRANSPORT startdma  ;
and2_1231: n_1524 <=  n_1525  AND n_1526;
delay_1232: n_1525  <= TRANSPORT a_LC1_C15  ;
delay_1233: n_1526  <= TRANSPORT startdma  ;
and1_1234: n_1527 <=  gnd;
delay_1235: n_1528  <= TRANSPORT clk  ;
filter_1236: FILTER_a8237

    PORT MAP (IN1 => n_1528, Y => a_N3553_aCLK);
dff_1237: DFF_a8237

    PORT MAP ( D => a_EQ1019, CLK => a_SCH2BAROUT_F8_G_aCLK, CLRN => a_SCH2BAROUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F8_G);
inv_1238: a_SCH2BAROUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1239: a_EQ1019 <=  n_1537  XOR n_1545;
or2_1240: n_1537 <=  n_1538  OR n_1542;
and2_1241: n_1538 <=  n_1539  AND n_1540;
inv_1242: n_1539  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_1243: n_1540  <= TRANSPORT dbin(0)  ;
and2_1244: n_1542 <=  n_1543  AND n_1544;
delay_1245: n_1543  <= TRANSPORT a_N2583_aNOT  ;
delay_1246: n_1544  <= TRANSPORT a_SCH2BAROUT_F8_G  ;
and1_1247: n_1545 <=  gnd;
delay_1248: n_1546  <= TRANSPORT clk  ;
filter_1249: FILTER_a8237

    PORT MAP (IN1 => n_1546, Y => a_SCH2BAROUT_F8_G_aCLK);
dff_1250: DFF_a8237

    PORT MAP ( D => a_EQ1099, CLK => a_SCH3BWORDOUT_F8_G_aCLK, CLRN => a_SCH3BWORDOUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F8_G);
inv_1251: a_SCH3BWORDOUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1252: a_EQ1099 <=  n_1555  XOR n_1562;
or2_1253: n_1555 <=  n_1556  OR n_1559;
and2_1254: n_1556 <=  n_1557  AND n_1558;
inv_1255: n_1557  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_1256: n_1558  <= TRANSPORT dbin(0)  ;
and2_1257: n_1559 <=  n_1560  AND n_1561;
delay_1258: n_1560  <= TRANSPORT a_N2573_aNOT  ;
delay_1259: n_1561  <= TRANSPORT a_SCH3BWORDOUT_F8_G  ;
and1_1260: n_1562 <=  gnd;
delay_1261: n_1563  <= TRANSPORT clk  ;
filter_1262: FILTER_a8237

    PORT MAP (IN1 => n_1563, Y => a_SCH3BWORDOUT_F8_G_aCLK);
delay_1263: a_N2354_aNOT  <= TRANSPORT a_N2354_aNOT_aIN  ;
xor2_1264: a_N2354_aNOT_aIN <=  n_1567  XOR n_1573;
or1_1265: n_1567 <=  n_1568;
and4_1266: n_1568 <=  n_1569  AND n_1570  AND n_1571  AND n_1572;
inv_1267: n_1569  <= TRANSPORT NOT ain(3)  ;
inv_1268: n_1570  <= TRANSPORT NOT ain(2)  ;
inv_1269: n_1571  <= TRANSPORT NOT ain(1)  ;
inv_1270: n_1572  <= TRANSPORT NOT ain(0)  ;
and1_1271: n_1573 <=  gnd;
delay_1272: a_N2586  <= TRANSPORT a_N2586_aIN  ;
xor2_1273: a_N2586_aIN <=  n_1576  XOR n_1581;
or1_1274: n_1576 <=  n_1577;
and2_1275: n_1577 <=  n_1578  AND n_1580;
inv_1276: n_1578  <= TRANSPORT NOT a_LC6_D6  ;
delay_1277: n_1580  <= TRANSPORT a_N2354_aNOT  ;
and1_1278: n_1581 <=  gnd;
delay_1279: a_N2587_aNOT  <= TRANSPORT a_EQ640  ;
xor2_1280: a_EQ640 <=  n_1584  XOR n_1589;
or2_1281: n_1584 <=  n_1585  OR n_1587;
and1_1282: n_1585 <=  n_1586;
inv_1283: n_1586  <= TRANSPORT NOT a_N2354_aNOT  ;
and1_1284: n_1587 <=  n_1588;
delay_1285: n_1588  <= TRANSPORT a_LC3_D22  ;
and1_1286: n_1589 <=  gnd;
dff_1287: DFF_a8237

    PORT MAP ( D => a_EQ891, CLK => a_SCH0BAROUT_F8_G_aCLK, CLRN => a_SCH0BAROUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F8_G);
inv_1288: a_SCH0BAROUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1289: a_EQ891 <=  n_1597  XOR n_1608;
or3_1290: n_1597 <=  n_1598  OR n_1602  OR n_1605;
and3_1291: n_1598 <=  n_1599  AND n_1600  AND n_1601;
inv_1292: n_1599  <= TRANSPORT NOT a_N2586  ;
inv_1293: n_1600  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_1294: n_1601  <= TRANSPORT dbin(0)  ;
and2_1295: n_1602 <=  n_1603  AND n_1604;
delay_1296: n_1603  <= TRANSPORT a_N2587_aNOT  ;
delay_1297: n_1604  <= TRANSPORT a_SCH0BAROUT_F8_G  ;
and2_1298: n_1605 <=  n_1606  AND n_1607;
delay_1299: n_1606  <= TRANSPORT a_N2586  ;
delay_1300: n_1607  <= TRANSPORT a_SCH0BAROUT_F8_G  ;
and1_1301: n_1608 <=  gnd;
delay_1302: n_1609  <= TRANSPORT clk  ;
filter_1303: FILTER_a8237

    PORT MAP (IN1 => n_1609, Y => a_SCH0BAROUT_F8_G_aCLK);
delay_1304: a_N2348  <= TRANSPORT a_EQ554  ;
xor2_1305: a_EQ554 <=  n_1613  XOR n_1622;
or4_1306: n_1613 <=  n_1614  OR n_1616  OR n_1618  OR n_1620;
and1_1307: n_1614 <=  n_1615;
delay_1308: n_1615  <= TRANSPORT ain(0)  ;
and1_1309: n_1616 <=  n_1617;
delay_1310: n_1617  <= TRANSPORT ain(3)  ;
and1_1311: n_1618 <=  n_1619;
inv_1312: n_1619  <= TRANSPORT NOT ain(2)  ;
and1_1313: n_1620 <=  n_1621;
inv_1314: n_1621  <= TRANSPORT NOT ain(1)  ;
and1_1315: n_1622 <=  gnd;
delay_1316: a_N2581_aNOT  <= TRANSPORT a_EQ632  ;
xor2_1317: a_EQ632 <=  n_1625  XOR n_1630;
or2_1318: n_1625 <=  n_1626  OR n_1628;
and1_1319: n_1626 <=  n_1627;
delay_1320: n_1627  <= TRANSPORT a_N2348  ;
and1_1321: n_1628 <=  n_1629;
delay_1322: n_1629  <= TRANSPORT a_LC3_D22  ;
and1_1323: n_1630 <=  gnd;
dff_1324: DFF_a8237

    PORT MAP ( D => a_EQ1083, CLK => a_SCH3BAROUT_F8_G_aCLK, CLRN => a_SCH3BAROUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F8_G);
inv_1325: a_SCH3BAROUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1326: a_EQ1083 <=  n_1638  XOR n_1645;
or2_1327: n_1638 <=  n_1639  OR n_1642;
and2_1328: n_1639 <=  n_1640  AND n_1641;
inv_1329: n_1640  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_1330: n_1641  <= TRANSPORT dbin(0)  ;
and2_1331: n_1642 <=  n_1643  AND n_1644;
delay_1332: n_1643  <= TRANSPORT a_N2581_aNOT  ;
delay_1333: n_1644  <= TRANSPORT a_SCH3BAROUT_F8_G  ;
and1_1334: n_1645 <=  gnd;
delay_1335: n_1646  <= TRANSPORT clk  ;
filter_1336: FILTER_a8237

    PORT MAP (IN1 => n_1646, Y => a_SCH3BAROUT_F8_G_aCLK);
dff_1337: DFF_a8237

    PORT MAP ( D => a_EQ907, CLK => a_SCH0BWORDOUT_F8_G_aCLK, CLRN => a_SCH0BWORDOUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F8_G);
inv_1338: a_SCH0BWORDOUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1339: a_EQ907 <=  n_1655  XOR n_1666;
or3_1340: n_1655 <=  n_1656  OR n_1660  OR n_1663;
and3_1341: n_1656 <=  n_1657  AND n_1658  AND n_1659;
inv_1342: n_1657  <= TRANSPORT NOT a_LC3_D22  ;
inv_1343: n_1658  <= TRANSPORT NOT a_N2353  ;
delay_1344: n_1659  <= TRANSPORT dbin(0)  ;
and2_1345: n_1660 <=  n_1661  AND n_1662;
delay_1346: n_1661  <= TRANSPORT a_N2353  ;
delay_1347: n_1662  <= TRANSPORT a_SCH0BWORDOUT_F8_G  ;
and2_1348: n_1663 <=  n_1664  AND n_1665;
delay_1349: n_1664  <= TRANSPORT a_LC3_D22  ;
delay_1350: n_1665  <= TRANSPORT a_SCH0BWORDOUT_F8_G  ;
and1_1351: n_1666 <=  gnd;
delay_1352: n_1667  <= TRANSPORT clk  ;
filter_1353: FILTER_a8237

    PORT MAP (IN1 => n_1667, Y => a_SCH0BWORDOUT_F8_G_aCLK);
dff_1354: DFF_a8237

    PORT MAP ( D => a_EQ955, CLK => a_SCH1BAROUT_F8_G_aCLK, CLRN => a_SCH1BAROUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F8_G);
inv_1355: a_SCH1BAROUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1356: a_EQ955 <=  n_1676  XOR n_1683;
or2_1357: n_1676 <=  n_1677  OR n_1680;
and2_1358: n_1677 <=  n_1678  AND n_1679;
inv_1359: n_1678  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_1360: n_1679  <= TRANSPORT dbin(0)  ;
and2_1361: n_1680 <=  n_1681  AND n_1682;
delay_1362: n_1681  <= TRANSPORT a_N2585_aNOT  ;
delay_1363: n_1682  <= TRANSPORT a_SCH1BAROUT_F8_G  ;
and1_1364: n_1683 <=  gnd;
delay_1365: n_1684  <= TRANSPORT clk  ;
filter_1366: FILTER_a8237

    PORT MAP (IN1 => n_1684, Y => a_SCH1BAROUT_F8_G_aCLK);
dff_1367: DFF_a8237

    PORT MAP ( D => a_EQ1035, CLK => a_SCH2BWORDOUT_F8_G_aCLK, CLRN => a_SCH2BWORDOUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F8_G);
inv_1368: a_SCH2BWORDOUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1369: a_EQ1035 <=  n_1693  XOR n_1704;
or3_1370: n_1693 <=  n_1694  OR n_1698  OR n_1701;
and3_1371: n_1694 <=  n_1695  AND n_1696  AND n_1697;
inv_1372: n_1695  <= TRANSPORT NOT a_LC3_D22  ;
inv_1373: n_1696  <= TRANSPORT NOT a_N62_aNOT  ;
delay_1374: n_1697  <= TRANSPORT dbin(0)  ;
and2_1375: n_1698 <=  n_1699  AND n_1700;
delay_1376: n_1699  <= TRANSPORT a_N62_aNOT  ;
delay_1377: n_1700  <= TRANSPORT a_SCH2BWORDOUT_F8_G  ;
and2_1378: n_1701 <=  n_1702  AND n_1703;
delay_1379: n_1702  <= TRANSPORT a_LC3_D22  ;
delay_1380: n_1703  <= TRANSPORT a_SCH2BWORDOUT_F8_G  ;
and1_1381: n_1704 <=  gnd;
delay_1382: n_1705  <= TRANSPORT clk  ;
filter_1383: FILTER_a8237

    PORT MAP (IN1 => n_1705, Y => a_SCH2BWORDOUT_F8_G_aCLK);
dff_1384: DFF_a8237

    PORT MAP ( D => a_EQ971, CLK => a_SCH1BWORDOUT_F8_G_aCLK, CLRN => a_SCH1BWORDOUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F8_G);
inv_1385: a_SCH1BWORDOUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1386: a_EQ971 <=  n_1714  XOR n_1721;
or2_1387: n_1714 <=  n_1715  OR n_1718;
and2_1388: n_1715 <=  n_1716  AND n_1717;
inv_1389: n_1716  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_1390: n_1717  <= TRANSPORT dbin(0)  ;
and2_1391: n_1718 <=  n_1719  AND n_1720;
delay_1392: n_1719  <= TRANSPORT a_N2577_aNOT  ;
delay_1393: n_1720  <= TRANSPORT a_SCH1BWORDOUT_F8_G  ;
and1_1394: n_1721 <=  gnd;
delay_1395: n_1722  <= TRANSPORT clk  ;
filter_1396: FILTER_a8237

    PORT MAP (IN1 => n_1722, Y => a_SCH1BWORDOUT_F8_G_aCLK);
dff_1397: DFF_a8237

    PORT MAP ( D => a_EQ1091, CLK => a_SCH3BWORDOUT_F0_G_aCLK, CLRN => a_SCH3BWORDOUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F0_G);
inv_1398: a_SCH3BWORDOUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1399: a_EQ1091 <=  n_1731  XOR n_1738;
or2_1400: n_1731 <=  n_1732  OR n_1735;
and2_1401: n_1732 <=  n_1733  AND n_1734;
inv_1402: n_1733  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_1403: n_1734  <= TRANSPORT dbin(0)  ;
and2_1404: n_1735 <=  n_1736  AND n_1737;
delay_1405: n_1736  <= TRANSPORT a_N2572_aNOT  ;
delay_1406: n_1737  <= TRANSPORT a_SCH3BWORDOUT_F0_G  ;
and1_1407: n_1738 <=  gnd;
delay_1408: n_1739  <= TRANSPORT clk  ;
filter_1409: FILTER_a8237

    PORT MAP (IN1 => n_1739, Y => a_SCH3BWORDOUT_F0_G_aCLK);
dff_1410: DFF_a8237

    PORT MAP ( D => a_EQ899, CLK => a_SCH0BWORDOUT_F0_G_aCLK, CLRN => a_SCH0BWORDOUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F0_G);
inv_1411: a_SCH0BWORDOUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1412: a_EQ899 <=  n_1748  XOR n_1755;
or2_1413: n_1748 <=  n_1749  OR n_1752;
and2_1414: n_1749 <=  n_1750  AND n_1751;
inv_1415: n_1750  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_1416: n_1751  <= TRANSPORT dbin(0)  ;
and2_1417: n_1752 <=  n_1753  AND n_1754;
delay_1418: n_1753  <= TRANSPORT a_N2578_aNOT  ;
delay_1419: n_1754  <= TRANSPORT a_SCH0BWORDOUT_F0_G  ;
and1_1420: n_1755 <=  gnd;
delay_1421: n_1756  <= TRANSPORT clk  ;
filter_1422: FILTER_a8237

    PORT MAP (IN1 => n_1756, Y => a_SCH0BWORDOUT_F0_G_aCLK);
dff_1423: DFF_a8237

    PORT MAP ( D => a_EQ1027, CLK => a_SCH2BWORDOUT_F0_G_aCLK, CLRN => a_SCH2BWORDOUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F0_G);
inv_1424: a_SCH2BWORDOUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1425: a_EQ1027 <=  n_1765  XOR n_1772;
or2_1426: n_1765 <=  n_1766  OR n_1769;
and2_1427: n_1766 <=  n_1767  AND n_1768;
inv_1428: n_1767  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_1429: n_1768  <= TRANSPORT dbin(0)  ;
and2_1430: n_1769 <=  n_1770  AND n_1771;
delay_1431: n_1770  <= TRANSPORT a_N2574_aNOT  ;
delay_1432: n_1771  <= TRANSPORT a_SCH2BWORDOUT_F0_G  ;
and1_1433: n_1772 <=  gnd;
delay_1434: n_1773  <= TRANSPORT clk  ;
filter_1435: FILTER_a8237

    PORT MAP (IN1 => n_1773, Y => a_SCH2BWORDOUT_F0_G_aCLK);
delay_1436: a_LC8_D12  <= TRANSPORT a_EQ516  ;
xor2_1437: a_EQ516 <=  n_1777  XOR n_1786;
or2_1438: n_1777 <=  n_1778  OR n_1782;
and2_1439: n_1778 <=  n_1779  AND n_1780;
inv_1440: n_1779  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_1441: n_1780  <= TRANSPORT a_SCH0WRDCNTREG_F0_G  ;
and2_1442: n_1782 <=  n_1783  AND n_1784;
delay_1443: n_1783  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_1444: n_1784  <= TRANSPORT a_SCH1WRDCNTREG_F0_G  ;
and1_1445: n_1786 <=  gnd;
delay_1446: a_N1867_aNOT  <= TRANSPORT a_EQ515  ;
xor2_1447: a_EQ515 <=  n_1789  XOR n_1801;
or3_1448: n_1789 <=  n_1790  OR n_1793  OR n_1797;
and2_1449: n_1790 <=  n_1791  AND n_1792;
delay_1450: n_1791  <= TRANSPORT a_N2531  ;
delay_1451: n_1792  <= TRANSPORT a_LC8_D12  ;
and3_1452: n_1793 <=  n_1794  AND n_1795  AND n_1796;
delay_1453: n_1794  <= TRANSPORT a_N2557  ;
inv_1454: n_1795  <= TRANSPORT NOT a_N2531  ;
inv_1455: n_1796  <= TRANSPORT NOT a_N3556  ;
and3_1456: n_1797 <=  n_1798  AND n_1799  AND n_1800;
inv_1457: n_1798  <= TRANSPORT NOT a_N2557  ;
inv_1458: n_1799  <= TRANSPORT NOT a_N2531  ;
delay_1459: n_1800  <= TRANSPORT a_N3556  ;
and1_1460: n_1801 <=  gnd;
delay_1461: a_LC5_D12  <= TRANSPORT a_EQ514  ;
xor2_1462: a_EQ514 <=  n_1804  XOR n_1812;
or2_1463: n_1804 <=  n_1805  OR n_1809;
and2_1464: n_1805 <=  n_1806  AND n_1807;
inv_1465: n_1806  <= TRANSPORT NOT a_N2377  ;
delay_1466: n_1807  <= TRANSPORT a_SCH3WRDCNTREG_F0_G  ;
and2_1467: n_1809 <=  n_1810  AND n_1811;
inv_1468: n_1810  <= TRANSPORT NOT a_N88_aNOT  ;
delay_1469: n_1811  <= TRANSPORT a_SCH1WRDCNTREG_F0_G  ;
and1_1470: n_1812 <=  gnd;
delay_1471: a_LC6_D12  <= TRANSPORT a_EQ513  ;
xor2_1472: a_EQ513 <=  n_1815  XOR n_1823;
or2_1473: n_1815 <=  n_1816  OR n_1819;
and2_1474: n_1816 <=  n_1817  AND n_1818;
inv_1475: n_1817  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_1476: n_1818  <= TRANSPORT a_SCH0WRDCNTREG_F0_G  ;
and2_1477: n_1819 <=  n_1820  AND n_1821;
inv_1478: n_1820  <= TRANSPORT NOT a_N2376  ;
delay_1479: n_1821  <= TRANSPORT a_SCH2WRDCNTREG_F0_G  ;
and1_1480: n_1823 <=  gnd;
dff_1481: DFF_a8237

    PORT MAP ( D => a_EQ852, CLK => a_N3556_aCLK, CLRN => a_N3556_aCLRN, PRN => vcc,
          Q => a_N3556);
inv_1482: a_N3556_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1483: a_EQ852 <=  n_1830  XOR n_1840;
or3_1484: n_1830 <=  n_1831  OR n_1834  OR n_1837;
and2_1485: n_1831 <=  n_1832  AND n_1833;
delay_1486: n_1832  <= TRANSPORT a_N1867_aNOT  ;
inv_1487: n_1833  <= TRANSPORT NOT startdma  ;
and2_1488: n_1834 <=  n_1835  AND n_1836;
delay_1489: n_1835  <= TRANSPORT a_LC5_D12  ;
delay_1490: n_1836  <= TRANSPORT startdma  ;
and2_1491: n_1837 <=  n_1838  AND n_1839;
delay_1492: n_1838  <= TRANSPORT a_LC6_D12  ;
delay_1493: n_1839  <= TRANSPORT startdma  ;
and1_1494: n_1840 <=  gnd;
delay_1495: n_1841  <= TRANSPORT clk  ;
filter_1496: FILTER_a8237

    PORT MAP (IN1 => n_1841, Y => a_N3556_aCLK);
dff_1497: DFF_a8237

    PORT MAP ( D => a_EQ1084, CLK => a_SCH3BAROUT_F9_G_aCLK, CLRN => a_SCH3BAROUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F9_G);
inv_1498: a_SCH3BAROUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1499: a_EQ1084 <=  n_1850  XOR n_1858;
or2_1500: n_1850 <=  n_1851  OR n_1855;
and2_1501: n_1851 <=  n_1852  AND n_1853;
inv_1502: n_1852  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_1503: n_1853  <= TRANSPORT dbin(1)  ;
and2_1504: n_1855 <=  n_1856  AND n_1857;
delay_1505: n_1856  <= TRANSPORT a_N2581_aNOT  ;
delay_1506: n_1857  <= TRANSPORT a_SCH3BAROUT_F9_G  ;
and1_1507: n_1858 <=  gnd;
delay_1508: n_1859  <= TRANSPORT clk  ;
filter_1509: FILTER_a8237

    PORT MAP (IN1 => n_1859, Y => a_SCH3BAROUT_F9_G_aCLK);
dff_1510: DFF_a8237

    PORT MAP ( D => a_EQ1020, CLK => a_SCH2BAROUT_F9_G_aCLK, CLRN => a_SCH2BAROUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F9_G);
inv_1511: a_SCH2BAROUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1512: a_EQ1020 <=  n_1868  XOR n_1875;
or2_1513: n_1868 <=  n_1869  OR n_1872;
and2_1514: n_1869 <=  n_1870  AND n_1871;
inv_1515: n_1870  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_1516: n_1871  <= TRANSPORT dbin(1)  ;
and2_1517: n_1872 <=  n_1873  AND n_1874;
delay_1518: n_1873  <= TRANSPORT a_N2583_aNOT  ;
delay_1519: n_1874  <= TRANSPORT a_SCH2BAROUT_F9_G  ;
and1_1520: n_1875 <=  gnd;
delay_1521: n_1876  <= TRANSPORT clk  ;
filter_1522: FILTER_a8237

    PORT MAP (IN1 => n_1876, Y => a_SCH2BAROUT_F9_G_aCLK);
dff_1523: DFF_a8237

    PORT MAP ( D => a_EQ892, CLK => a_SCH0BAROUT_F9_G_aCLK, CLRN => a_SCH0BAROUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F9_G);
inv_1524: a_SCH0BAROUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1525: a_EQ892 <=  n_1885  XOR n_1892;
or2_1526: n_1885 <=  n_1886  OR n_1889;
and2_1527: n_1886 <=  n_1887  AND n_1888;
inv_1528: n_1887  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_1529: n_1888  <= TRANSPORT dbin(1)  ;
and2_1530: n_1889 <=  n_1890  AND n_1891;
delay_1531: n_1890  <= TRANSPORT a_N2587_aNOT  ;
delay_1532: n_1891  <= TRANSPORT a_SCH0BAROUT_F9_G  ;
and1_1533: n_1892 <=  gnd;
delay_1534: n_1893  <= TRANSPORT clk  ;
filter_1535: FILTER_a8237

    PORT MAP (IN1 => n_1893, Y => a_SCH0BAROUT_F9_G_aCLK);
delay_1536: a_LC3_C13  <= TRANSPORT a_EQ036  ;
xor2_1537: a_EQ036 <=  n_1897  XOR n_1906;
or4_1538: n_1897 <=  n_1898  OR n_1900  OR n_1902  OR n_1904;
and1_1539: n_1898 <=  n_1899;
delay_1540: n_1899  <= TRANSPORT a_N3554  ;
and1_1541: n_1900 <=  n_1901;
delay_1542: n_1901  <= TRANSPORT a_N3556  ;
and1_1543: n_1902 <=  n_1903;
delay_1544: n_1903  <= TRANSPORT a_N3555  ;
and1_1545: n_1904 <=  n_1905;
delay_1546: n_1905  <= TRANSPORT a_N3553  ;
and1_1547: n_1906 <=  gnd;
delay_1548: a_LC8_F13_aNOT  <= TRANSPORT a_LC8_F13_aNOT_aIN  ;
xor2_1549: a_LC8_F13_aNOT_aIN <=  n_1909  XOR n_1918;
or1_1550: n_1909 <=  n_1910;
and4_1551: n_1910 <=  n_1911  AND n_1912  AND n_1914  AND n_1916;
inv_1552: n_1911  <= TRANSPORT NOT a_LC3_C13  ;
inv_1553: n_1912  <= TRANSPORT NOT a_N3552  ;
inv_1554: n_1914  <= TRANSPORT NOT a_N3551  ;
inv_1555: n_1916  <= TRANSPORT NOT a_N3550  ;
and1_1556: n_1918 <=  gnd;
delay_1557: a_LC4_A13_aNOT  <= TRANSPORT a_LC4_A13_aNOT_aIN  ;
xor2_1558: a_LC4_A13_aNOT_aIN <=  n_1921  XOR n_1930;
or1_1559: n_1921 <=  n_1922;
and4_1560: n_1922 <=  n_1923  AND n_1924  AND n_1926  AND n_1928;
delay_1561: n_1923  <= TRANSPORT a_LC8_F13_aNOT  ;
inv_1562: n_1924  <= TRANSPORT NOT a_N3549  ;
inv_1563: n_1926  <= TRANSPORT NOT a_N3548  ;
inv_1564: n_1928  <= TRANSPORT NOT a_N3547  ;
and1_1565: n_1930 <=  gnd;
delay_1566: a_LC1_A20_aNOT  <= TRANSPORT a_LC1_A20_aNOT_aIN  ;
xor2_1567: a_LC1_A20_aNOT_aIN <=  n_1933  XOR n_1942;
or1_1568: n_1933 <=  n_1934;
and4_1569: n_1934 <=  n_1935  AND n_1936  AND n_1938  AND n_1940;
delay_1570: n_1935  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_1571: n_1936  <= TRANSPORT NOT a_N3546  ;
inv_1572: n_1938  <= TRANSPORT NOT a_N3545  ;
inv_1573: n_1940  <= TRANSPORT NOT a_N3544  ;
and1_1574: n_1942 <=  gnd;
delay_1575: a_LC3_E16_aNOT  <= TRANSPORT a_LC3_E16_aNOT_aIN  ;
xor2_1576: a_LC3_E16_aNOT_aIN <=  n_1945  XOR n_1952;
or1_1577: n_1945 <=  n_1946;
and3_1578: n_1946 <=  n_1947  AND n_1948  AND n_1950;
delay_1579: n_1947  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_1580: n_1948  <= TRANSPORT NOT a_N3543  ;
inv_1581: n_1950  <= TRANSPORT NOT a_N3542  ;
and1_1582: n_1952 <=  gnd;
delay_1583: a_N2539  <= TRANSPORT a_N2539_aIN  ;
xor2_1584: a_N2539_aIN <=  n_1955  XOR n_1960;
or1_1585: n_1955 <=  n_1956;
and2_1586: n_1956 <=  n_1957  AND n_1958;
delay_1587: n_1957  <= TRANSPORT a_LC3_E16_aNOT  ;
inv_1588: n_1958  <= TRANSPORT NOT a_N3541  ;
and1_1589: n_1960 <=  gnd;
delay_1590: a_LC1_B12  <= TRANSPORT a_EQ1164  ;
xor2_1591: a_EQ1164 <=  n_1963  XOR n_1980;
or4_1592: n_1963 <=  n_1964  OR n_1968  OR n_1972  OR n_1976;
and3_1593: n_1964 <=  n_1965  AND n_1966  AND n_1967;
inv_1594: n_1965  <= TRANSPORT NOT a_N820  ;
delay_1595: n_1966  <= TRANSPORT a_N822  ;
inv_1596: n_1967  <= TRANSPORT NOT a_N823  ;
and3_1597: n_1968 <=  n_1969  AND n_1970  AND n_1971;
inv_1598: n_1969  <= TRANSPORT NOT a_N820  ;
inv_1599: n_1970  <= TRANSPORT NOT a_N822  ;
inv_1600: n_1971  <= TRANSPORT NOT a_N821  ;
and3_1601: n_1972 <=  n_1973  AND n_1974  AND n_1975;
delay_1602: n_1973  <= TRANSPORT a_N820  ;
delay_1603: n_1974  <= TRANSPORT a_N821  ;
inv_1604: n_1975  <= TRANSPORT NOT a_N823  ;
and3_1605: n_1976 <=  n_1977  AND n_1978  AND n_1979;
delay_1606: n_1977  <= TRANSPORT a_N820  ;
inv_1607: n_1978  <= TRANSPORT NOT a_N822  ;
delay_1608: n_1979  <= TRANSPORT a_N821  ;
and1_1609: n_1980 <=  gnd;
delay_1610: a_SNEOPOUT_aNOT  <= TRANSPORT a_EQ1163  ;
xor2_1611: a_EQ1163 <=  n_1982  XOR n_1991;
or2_1612: n_1982 <=  n_1983  OR n_1987;
and3_1613: n_1983 <=  n_1984  AND n_1985  AND n_1986;
delay_1614: n_1984  <= TRANSPORT a_N1588  ;
delay_1615: n_1985  <= TRANSPORT a_N2539  ;
delay_1616: n_1986  <= TRANSPORT a_LC1_B12  ;
and3_1617: n_1987 <=  n_1988  AND n_1989  AND n_1990;
delay_1618: n_1988  <= TRANSPORT a_LC1_B23_aNOT  ;
delay_1619: n_1989  <= TRANSPORT a_N1588  ;
delay_1620: n_1990  <= TRANSPORT a_LC1_B12  ;
and1_1621: n_1991 <=  gnd;
delay_1622: a_N57_aNOT  <= TRANSPORT a_EQ181  ;
xor2_1623: a_EQ181 <=  n_1994  XOR n_2001;
or2_1624: n_1994 <=  n_1995  OR n_1997;
and1_1625: n_1995 <=  n_1996;
delay_1626: n_1996  <= TRANSPORT a_SNEOPOUT_aNOT  ;
and2_1627: n_1997 <=  n_1998  AND n_1999;
inv_1628: n_1998  <= TRANSPORT NOT a_LC1_B23_aNOT  ;
delay_1629: n_1999  <= TRANSPORT a_N825  ;
and1_1630: n_2001 <=  gnd;
delay_1631: a_N2528  <= TRANSPORT a_N2528_aIN  ;
xor2_1632: a_N2528_aIN <=  n_2004  XOR n_2009;
or1_1633: n_2004 <=  n_2005;
and2_1634: n_2005 <=  n_2006  AND n_2007;
delay_1635: n_2006  <= TRANSPORT a_N57_aNOT  ;
delay_1636: n_2007  <= TRANSPORT a_SCH3MODEREG_F2_G  ;
and1_1637: n_2009 <=  gnd;
delay_1638: a_N965  <= TRANSPORT a_EQ331  ;
xor2_1639: a_EQ331 <=  n_2012  XOR n_2017;
or2_1640: n_2012 <=  n_2013  OR n_2015;
and1_1641: n_2013 <=  n_2014;
inv_1642: n_2014  <= TRANSPORT NOT a_N2557  ;
and1_1643: n_2015 <=  n_2016;
delay_1644: n_2016  <= TRANSPORT a_N2377  ;
and1_1645: n_2017 <=  gnd;
delay_1646: a_N1095  <= TRANSPORT a_N1095_aIN  ;
xor2_1647: a_N1095_aIN <=  n_2020  XOR n_2024;
or1_1648: n_2020 <=  n_2021;
and2_1649: n_2021 <=  n_2022  AND n_2023;
inv_1650: n_2022  <= TRANSPORT NOT a_N2528  ;
delay_1651: n_2023  <= TRANSPORT a_N965  ;
and1_1652: n_2024 <=  gnd;
delay_1653: a_LC3_C4  <= TRANSPORT a_EQ832  ;
xor2_1654: a_EQ832 <=  n_2027  XOR n_2036;
or2_1655: n_2027 <=  n_2028  OR n_2032;
and3_1656: n_2028 <=  n_2029  AND n_2030  AND n_2031;
inv_1657: n_2029  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_1658: n_2030  <= TRANSPORT a_N1095  ;
delay_1659: n_2031  <= TRANSPORT dbin(1)  ;
and3_1660: n_2032 <=  n_2033  AND n_2034  AND n_2035;
delay_1661: n_2033  <= TRANSPORT a_N2572_aNOT  ;
delay_1662: n_2034  <= TRANSPORT a_N1095  ;
delay_1663: n_2035  <= TRANSPORT a_SCH3WRDCNTREG_F1_G  ;
and1_1664: n_2036 <=  gnd;
delay_1665: a_N1046_aNOT  <= TRANSPORT a_N1046_aNOT_aIN  ;
xor2_1666: a_N1046_aNOT_aIN <=  n_2039  XOR n_2044;
or1_1667: n_2039 <=  n_2040;
and2_1668: n_2040 <=  n_2041  AND n_2043;
delay_1669: n_2041  <= TRANSPORT a_SCH3BWORDOUT_F1_G  ;
delay_1670: n_2043  <= TRANSPORT a_N2528  ;
and1_1671: n_2044 <=  gnd;
delay_1672: a_N1094  <= TRANSPORT a_N1094_aIN  ;
xor2_1673: a_N1094_aIN <=  n_2047  XOR n_2051;
or1_1674: n_2047 <=  n_2048;
and2_1675: n_2048 <=  n_2049  AND n_2050;
inv_1676: n_2049  <= TRANSPORT NOT a_N2528  ;
inv_1677: n_2050  <= TRANSPORT NOT a_N965  ;
and1_1678: n_2051 <=  gnd;
dff_1679: DFF_a8237

    PORT MAP ( D => a_EQ1114, CLK => a_SCH3WRDCNTREG_F1_G_aCLK, CLRN => a_SCH3WRDCNTREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F1_G);
inv_1680: a_SCH3WRDCNTREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1681: a_EQ1114 <=  n_2058  XOR n_2066;
or3_1682: n_2058 <=  n_2059  OR n_2061  OR n_2063;
and1_1683: n_2059 <=  n_2060;
delay_1684: n_2060  <= TRANSPORT a_LC3_C4  ;
and1_1685: n_2061 <=  n_2062;
delay_1686: n_2062  <= TRANSPORT a_N1046_aNOT  ;
and2_1687: n_2063 <=  n_2064  AND n_2065;
inv_1688: n_2064  <= TRANSPORT NOT a_LC7_C22  ;
delay_1689: n_2065  <= TRANSPORT a_N1094  ;
and1_1690: n_2066 <=  gnd;
delay_1691: n_2067  <= TRANSPORT clk  ;
filter_1692: FILTER_a8237

    PORT MAP (IN1 => n_2067, Y => a_SCH3WRDCNTREG_F1_G_aCLK);
delay_1693: a_N2558_aNOT  <= TRANSPORT a_EQ613  ;
xor2_1694: a_EQ613 <=  n_2071  XOR n_2079;
or3_1695: n_2071 <=  n_2072  OR n_2075  OR n_2077;
and2_1696: n_2072 <=  n_2073  AND n_2074;
inv_1697: n_2073  <= TRANSPORT NOT a_N71_aNOT  ;
delay_1698: n_2074  <= TRANSPORT a_N2591  ;
and1_1699: n_2075 <=  n_2076;
delay_1700: n_2076  <= TRANSPORT a_N2598_aNOT  ;
and1_1701: n_2077 <=  n_2078;
inv_1702: n_2078  <= TRANSPORT NOT a_N2557  ;
and1_1703: n_2079 <=  gnd;
delay_1704: a_LC1_C12  <= TRANSPORT a_EQ771  ;
xor2_1705: a_EQ771 <=  n_2082  XOR n_2093;
or3_1706: n_2082 <=  n_2083  OR n_2087  OR n_2090;
and3_1707: n_2083 <=  n_2084  AND n_2085  AND n_2086;
inv_1708: n_2084  <= TRANSPORT NOT a_LC6_D6  ;
inv_1709: n_2085  <= TRANSPORT NOT a_N2353  ;
delay_1710: n_2086  <= TRANSPORT dbin(1)  ;
and2_1711: n_2087 <=  n_2088  AND n_2089;
delay_1712: n_2088  <= TRANSPORT a_N2353  ;
delay_1713: n_2089  <= TRANSPORT a_SCH0WRDCNTREG_F1_G  ;
and2_1714: n_2090 <=  n_2091  AND n_2092;
delay_1715: n_2091  <= TRANSPORT a_LC6_D6  ;
delay_1716: n_2092  <= TRANSPORT a_SCH0WRDCNTREG_F1_G  ;
and1_1717: n_2093 <=  gnd;
delay_1718: a_LC2_C12  <= TRANSPORT a_EQ772  ;
xor2_1719: a_EQ772 <=  n_2096  XOR n_2103;
or2_1720: n_2096 <=  n_2097  OR n_2100;
and2_1721: n_2097 <=  n_2098  AND n_2099;
inv_1722: n_2098  <= TRANSPORT NOT a_LC7_C22  ;
inv_1723: n_2099  <= TRANSPORT NOT a_N2558_aNOT  ;
and2_1724: n_2100 <=  n_2101  AND n_2102;
delay_1725: n_2101  <= TRANSPORT a_N2558_aNOT  ;
delay_1726: n_2102  <= TRANSPORT a_LC1_C12  ;
and1_1727: n_2103 <=  gnd;
delay_1728: a_N2525  <= TRANSPORT a_N2525_aIN  ;
xor2_1729: a_N2525_aIN <=  n_2106  XOR n_2111;
or1_1730: n_2106 <=  n_2107;
and2_1731: n_2107 <=  n_2108  AND n_2109;
delay_1732: n_2108  <= TRANSPORT a_N57_aNOT  ;
delay_1733: n_2109  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and1_1734: n_2111 <=  gnd;
dff_1735: DFF_a8237

    PORT MAP ( D => a_EQ922, CLK => a_SCH0WRDCNTREG_F1_G_aCLK, CLRN => a_SCH0WRDCNTREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F1_G);
inv_1736: a_SCH0WRDCNTREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1737: a_EQ922 <=  n_2118  XOR n_2126;
or2_1738: n_2118 <=  n_2119  OR n_2122;
and2_1739: n_2119 <=  n_2120  AND n_2121;
delay_1740: n_2120  <= TRANSPORT a_LC2_C12  ;
inv_1741: n_2121  <= TRANSPORT NOT a_N2525  ;
and2_1742: n_2122 <=  n_2123  AND n_2125;
delay_1743: n_2123  <= TRANSPORT a_SCH0BWORDOUT_F1_G  ;
delay_1744: n_2125  <= TRANSPORT a_N2525  ;
and1_1745: n_2126 <=  gnd;
delay_1746: n_2127  <= TRANSPORT clk  ;
filter_1747: FILTER_a8237

    PORT MAP (IN1 => n_2127, Y => a_SCH0WRDCNTREG_F1_G_aCLK);
delay_1748: a_N2559_aNOT  <= TRANSPORT a_EQ614  ;
xor2_1749: a_EQ614 <=  n_2131  XOR n_2140;
or3_1750: n_2131 <=  n_2132  OR n_2135  OR n_2138;
and2_1751: n_2132 <=  n_2133  AND n_2134;
inv_1752: n_2133  <= TRANSPORT NOT a_N2591  ;
delay_1753: n_2134  <= TRANSPORT a_N88_aNOT  ;
and2_1754: n_2135 <=  n_2136  AND n_2137;
delay_1755: n_2136  <= TRANSPORT a_N71_aNOT  ;
delay_1756: n_2137  <= TRANSPORT a_N88_aNOT  ;
and1_1757: n_2138 <=  n_2139;
inv_1758: n_2139  <= TRANSPORT NOT a_N2557  ;
and1_1759: n_2140 <=  gnd;
delay_1760: a_N2526  <= TRANSPORT a_N2526_aIN  ;
xor2_1761: a_N2526_aIN <=  n_2143  XOR n_2148;
or1_1762: n_2143 <=  n_2144;
and2_1763: n_2144 <=  n_2145  AND n_2146;
delay_1764: n_2145  <= TRANSPORT a_N57_aNOT  ;
delay_1765: n_2146  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and1_1766: n_2148 <=  gnd;
delay_1767: a_N2595  <= TRANSPORT a_N2595_aIN  ;
xor2_1768: a_N2595_aIN <=  n_2151  XOR n_2155;
or1_1769: n_2151 <=  n_2152;
and2_1770: n_2152 <=  n_2153  AND n_2154;
delay_1771: n_2153  <= TRANSPORT a_N2559_aNOT  ;
inv_1772: n_2154  <= TRANSPORT NOT a_N2526  ;
and1_1773: n_2155 <=  gnd;
delay_1774: a_LC7_D26  <= TRANSPORT a_LC7_D26_aIN  ;
xor2_1775: a_LC7_D26_aIN <=  n_2158  XOR n_2162;
or1_1776: n_2158 <=  n_2159;
and2_1777: n_2159 <=  n_2160  AND n_2161;
delay_1778: n_2160  <= TRANSPORT a_N2576_aNOT  ;
delay_1779: n_2161  <= TRANSPORT a_N2595  ;
and1_1780: n_2162 <=  gnd;
delay_1781: a_LC6_A25  <= TRANSPORT a_EQ793  ;
xor2_1782: a_EQ793 <=  n_2165  XOR n_2173;
or2_1783: n_2165 <=  n_2166  OR n_2169;
and2_1784: n_2166 <=  n_2167  AND n_2168;
delay_1785: n_2167  <= TRANSPORT a_LC7_D26  ;
delay_1786: n_2168  <= TRANSPORT a_SCH1WRDCNTREG_F1_G  ;
and2_1787: n_2169 <=  n_2170  AND n_2172;
delay_1788: n_2170  <= TRANSPORT a_SCH1BWORDOUT_F1_G  ;
delay_1789: n_2172  <= TRANSPORT a_N2526  ;
and1_1790: n_2173 <=  gnd;
delay_1791: a_N433  <= TRANSPORT a_N433_aIN  ;
xor2_1792: a_N433_aIN <=  n_2176  XOR n_2182;
or1_1793: n_2176 <=  n_2177;
and4_1794: n_2177 <=  n_2178  AND n_2179  AND n_2180  AND n_2181;
inv_1795: n_2178  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_1796: n_2179  <= TRANSPORT a_N2559_aNOT  ;
inv_1797: n_2180  <= TRANSPORT NOT a_N2526  ;
delay_1798: n_2181  <= TRANSPORT dbin(1)  ;
and1_1799: n_2182 <=  gnd;
delay_1800: a_N460  <= TRANSPORT a_N460_aIN  ;
xor2_1801: a_N460_aIN <=  n_2185  XOR n_2189;
or1_1802: n_2185 <=  n_2186;
and2_1803: n_2186 <=  n_2187  AND n_2188;
inv_1804: n_2187  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_1805: n_2188  <= TRANSPORT NOT a_N2526  ;
and1_1806: n_2189 <=  gnd;
dff_1807: DFF_a8237

    PORT MAP ( D => a_EQ986, CLK => a_SCH1WRDCNTREG_F1_G_aCLK, CLRN => a_SCH1WRDCNTREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F1_G);
inv_1808: a_SCH1WRDCNTREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1809: a_EQ986 <=  n_2196  XOR n_2204;
or3_1810: n_2196 <=  n_2197  OR n_2199  OR n_2201;
and1_1811: n_2197 <=  n_2198;
delay_1812: n_2198  <= TRANSPORT a_LC6_A25  ;
and1_1813: n_2199 <=  n_2200;
delay_1814: n_2200  <= TRANSPORT a_N433  ;
and2_1815: n_2201 <=  n_2202  AND n_2203;
inv_1816: n_2202  <= TRANSPORT NOT a_LC7_C22  ;
delay_1817: n_2203  <= TRANSPORT a_N460  ;
and1_1818: n_2204 <=  gnd;
delay_1819: n_2205  <= TRANSPORT clk  ;
filter_1820: FILTER_a8237

    PORT MAP (IN1 => n_2205, Y => a_SCH1WRDCNTREG_F1_G_aCLK);
delay_1821: a_N2560_aNOT  <= TRANSPORT a_EQ615  ;
xor2_1822: a_EQ615 <=  n_2209  XOR n_2214;
or2_1823: n_2209 <=  n_2210  OR n_2212;
and1_1824: n_2210 <=  n_2211;
inv_1825: n_2211  <= TRANSPORT NOT a_N2557  ;
and1_1826: n_2212 <=  n_2213;
delay_1827: n_2213  <= TRANSPORT a_N2376  ;
and1_1828: n_2214 <=  gnd;
delay_1829: a_N2527  <= TRANSPORT a_N2527_aIN  ;
xor2_1830: a_N2527_aIN <=  n_2217  XOR n_2222;
or1_1831: n_2217 <=  n_2218;
and2_1832: n_2218 <=  n_2219  AND n_2220;
delay_1833: n_2219  <= TRANSPORT a_N57_aNOT  ;
delay_1834: n_2220  <= TRANSPORT a_SCH2MODEREG_F2_G  ;
and1_1835: n_2222 <=  gnd;
delay_1836: a_N756  <= TRANSPORT a_N756_aIN  ;
xor2_1837: a_N756_aIN <=  n_2225  XOR n_2229;
or1_1838: n_2225 <=  n_2226;
and2_1839: n_2226 <=  n_2227  AND n_2228;
delay_1840: n_2227  <= TRANSPORT a_N2560_aNOT  ;
inv_1841: n_2228  <= TRANSPORT NOT a_N2527  ;
and1_1842: n_2229 <=  gnd;
delay_1843: a_LC2_C18  <= TRANSPORT a_EQ812  ;
xor2_1844: a_EQ812 <=  n_2232  XOR n_2241;
or2_1845: n_2232 <=  n_2233  OR n_2237;
and3_1846: n_2233 <=  n_2234  AND n_2235  AND n_2236;
inv_1847: n_2234  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_1848: n_2235  <= TRANSPORT a_N756  ;
delay_1849: n_2236  <= TRANSPORT dbin(1)  ;
and3_1850: n_2237 <=  n_2238  AND n_2239  AND n_2240;
delay_1851: n_2238  <= TRANSPORT a_N2574_aNOT  ;
delay_1852: n_2239  <= TRANSPORT a_N756  ;
delay_1853: n_2240  <= TRANSPORT a_SCH2WRDCNTREG_F1_G  ;
and1_1854: n_2241 <=  gnd;
delay_1855: a_N797  <= TRANSPORT a_N797_aIN  ;
xor2_1856: a_N797_aIN <=  n_2244  XOR n_2249;
or1_1857: n_2244 <=  n_2245;
and2_1858: n_2245 <=  n_2246  AND n_2248;
delay_1859: n_2246  <= TRANSPORT a_SCH2BWORDOUT_F1_G  ;
delay_1860: n_2248  <= TRANSPORT a_N2527  ;
and1_1861: n_2249 <=  gnd;
delay_1862: a_N858  <= TRANSPORT a_N858_aIN  ;
xor2_1863: a_N858_aIN <=  n_2252  XOR n_2256;
or1_1864: n_2252 <=  n_2253;
and2_1865: n_2253 <=  n_2254  AND n_2255;
inv_1866: n_2254  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_1867: n_2255  <= TRANSPORT NOT a_N2527  ;
and1_1868: n_2256 <=  gnd;
dff_1869: DFF_a8237

    PORT MAP ( D => a_EQ1050, CLK => a_SCH2WRDCNTREG_F1_G_aCLK, CLRN => a_SCH2WRDCNTREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F1_G);
inv_1870: a_SCH2WRDCNTREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1871: a_EQ1050 <=  n_2263  XOR n_2271;
or3_1872: n_2263 <=  n_2264  OR n_2266  OR n_2268;
and1_1873: n_2264 <=  n_2265;
delay_1874: n_2265  <= TRANSPORT a_LC2_C18  ;
and1_1875: n_2266 <=  n_2267;
delay_1876: n_2267  <= TRANSPORT a_N797  ;
and2_1877: n_2268 <=  n_2269  AND n_2270;
inv_1878: n_2269  <= TRANSPORT NOT a_LC7_C22  ;
delay_1879: n_2270  <= TRANSPORT a_N858  ;
and1_1880: n_2271 <=  gnd;
delay_1881: n_2272  <= TRANSPORT clk  ;
filter_1882: FILTER_a8237

    PORT MAP (IN1 => n_2272, Y => a_SCH2WRDCNTREG_F1_G_aCLK);
delay_1883: a_LC1_A13  <= TRANSPORT a_EQ028  ;
xor2_1884: a_EQ028 <=  n_2276  XOR n_2291;
or4_1885: n_2276 <=  n_2277  OR n_2280  OR n_2283  OR n_2286;
and2_1886: n_2277 <=  n_2278  AND n_2279;
delay_1887: n_2278  <= TRANSPORT a_N3548  ;
inv_1888: n_2279  <= TRANSPORT NOT a_N3547  ;
and2_1889: n_2280 <=  n_2281  AND n_2282;
delay_1890: n_2281  <= TRANSPORT a_N3549  ;
inv_1891: n_2282  <= TRANSPORT NOT a_N3547  ;
and2_1892: n_2283 <=  n_2284  AND n_2285;
inv_1893: n_2284  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
inv_1894: n_2285  <= TRANSPORT NOT a_N3547  ;
and4_1895: n_2286 <=  n_2287  AND n_2288  AND n_2289  AND n_2290;
delay_1896: n_2287  <= TRANSPORT a_LC8_F13_aNOT  ;
inv_1897: n_2288  <= TRANSPORT NOT a_N3549  ;
inv_1898: n_2289  <= TRANSPORT NOT a_N3548  ;
delay_1899: n_2290  <= TRANSPORT a_N3547  ;
and1_1900: n_2291 <=  gnd;
delay_1901: a_LC3_A7  <= TRANSPORT a_EQ758  ;
xor2_1902: a_EQ758 <=  n_2294  XOR n_2306;
or3_1903: n_2294 <=  n_2295  OR n_2299  OR n_2303;
and3_1904: n_2295 <=  n_2296  AND n_2297  AND n_2298;
inv_1905: n_2296  <= TRANSPORT NOT a_LC3_D22  ;
inv_1906: n_2297  <= TRANSPORT NOT a_N2353  ;
delay_1907: n_2298  <= TRANSPORT dbin(1)  ;
and2_1908: n_2299 <=  n_2300  AND n_2301;
delay_1909: n_2300  <= TRANSPORT a_N2353  ;
delay_1910: n_2301  <= TRANSPORT a_SCH0WRDCNTREG_F9_G  ;
and2_1911: n_2303 <=  n_2304  AND n_2305;
delay_1912: n_2304  <= TRANSPORT a_LC3_D22  ;
delay_1913: n_2305  <= TRANSPORT a_SCH0WRDCNTREG_F9_G  ;
and1_1914: n_2306 <=  gnd;
delay_1915: a_LC4_A7  <= TRANSPORT a_EQ759  ;
xor2_1916: a_EQ759 <=  n_2309  XOR n_2316;
or2_1917: n_2309 <=  n_2310  OR n_2313;
and2_1918: n_2310 <=  n_2311  AND n_2312;
inv_1919: n_2311  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_1920: n_2312  <= TRANSPORT NOT a_LC1_A13  ;
and2_1921: n_2313 <=  n_2314  AND n_2315;
delay_1922: n_2314  <= TRANSPORT a_N2558_aNOT  ;
delay_1923: n_2315  <= TRANSPORT a_LC3_A7  ;
and1_1924: n_2316 <=  gnd;
dff_1925: DFF_a8237

    PORT MAP ( D => a_EQ930, CLK => a_SCH0WRDCNTREG_F9_G_aCLK, CLRN => a_SCH0WRDCNTREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F9_G);
inv_1926: a_SCH0WRDCNTREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1927: a_EQ930 <=  n_2323  XOR n_2331;
or2_1928: n_2323 <=  n_2324  OR n_2327;
and2_1929: n_2324 <=  n_2325  AND n_2326;
inv_1930: n_2325  <= TRANSPORT NOT a_N2525  ;
delay_1931: n_2326  <= TRANSPORT a_LC4_A7  ;
and2_1932: n_2327 <=  n_2328  AND n_2330;
delay_1933: n_2328  <= TRANSPORT a_SCH0BWORDOUT_F9_G  ;
delay_1934: n_2330  <= TRANSPORT a_N2525  ;
and1_1935: n_2331 <=  gnd;
delay_1936: n_2332  <= TRANSPORT clk  ;
filter_1937: FILTER_a8237

    PORT MAP (IN1 => n_2332, Y => a_SCH0WRDCNTREG_F9_G_aCLK);
delay_1938: a_LC2_E12  <= TRANSPORT a_LC2_E12_aIN  ;
xor2_1939: a_LC2_E12_aIN <=  n_2336  XOR n_2340;
or1_1940: n_2336 <=  n_2337;
and2_1941: n_2337 <=  n_2338  AND n_2339;
delay_1942: n_2338  <= TRANSPORT a_N2577_aNOT  ;
delay_1943: n_2339  <= TRANSPORT a_N2595  ;
and1_1944: n_2340 <=  gnd;
delay_1945: a_LC3_A25  <= TRANSPORT a_EQ782  ;
xor2_1946: a_EQ782 <=  n_2343  XOR n_2352;
or2_1947: n_2343 <=  n_2344  OR n_2348;
and2_1948: n_2344 <=  n_2345  AND n_2346;
delay_1949: n_2345  <= TRANSPORT a_LC2_E12  ;
delay_1950: n_2346  <= TRANSPORT a_SCH1WRDCNTREG_F9_G  ;
and2_1951: n_2348 <=  n_2349  AND n_2351;
delay_1952: n_2349  <= TRANSPORT a_SCH1BWORDOUT_F9_G  ;
delay_1953: n_2351  <= TRANSPORT a_N2526  ;
and1_1954: n_2352 <=  gnd;
delay_1955: a_N636_aNOT  <= TRANSPORT a_N636_aNOT_aIN  ;
xor2_1956: a_N636_aNOT_aIN <=  n_2355  XOR n_2361;
or1_1957: n_2355 <=  n_2356;
and4_1958: n_2356 <=  n_2357  AND n_2358  AND n_2359  AND n_2360;
inv_1959: n_2357  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_1960: n_2358  <= TRANSPORT a_N2559_aNOT  ;
inv_1961: n_2359  <= TRANSPORT NOT a_N2526  ;
delay_1962: n_2360  <= TRANSPORT dbin(1)  ;
and1_1963: n_2361 <=  gnd;
dff_1964: DFF_a8237

    PORT MAP ( D => a_EQ994, CLK => a_SCH1WRDCNTREG_F9_G_aCLK, CLRN => a_SCH1WRDCNTREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F9_G);
inv_1965: a_SCH1WRDCNTREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_1966: a_EQ994 <=  n_2368  XOR n_2376;
or3_1967: n_2368 <=  n_2369  OR n_2371  OR n_2373;
and1_1968: n_2369 <=  n_2370;
delay_1969: n_2370  <= TRANSPORT a_LC3_A25  ;
and1_1970: n_2371 <=  n_2372;
delay_1971: n_2372  <= TRANSPORT a_N636_aNOT  ;
and2_1972: n_2373 <=  n_2374  AND n_2375;
delay_1973: n_2374  <= TRANSPORT a_N460  ;
inv_1974: n_2375  <= TRANSPORT NOT a_LC1_A13  ;
and1_1975: n_2376 <=  gnd;
delay_1976: n_2377  <= TRANSPORT clk  ;
filter_1977: FILTER_a8237

    PORT MAP (IN1 => n_2377, Y => a_SCH1WRDCNTREG_F9_G_aCLK);
delay_1978: a_LC1_A7  <= TRANSPORT a_EQ803  ;
xor2_1979: a_EQ803 <=  n_2381  XOR n_2393;
or3_1980: n_2381 <=  n_2382  OR n_2386  OR n_2390;
and3_1981: n_2382 <=  n_2383  AND n_2384  AND n_2385;
inv_1982: n_2383  <= TRANSPORT NOT a_LC3_D22  ;
inv_1983: n_2384  <= TRANSPORT NOT a_N62_aNOT  ;
delay_1984: n_2385  <= TRANSPORT dbin(1)  ;
and2_1985: n_2386 <=  n_2387  AND n_2388;
delay_1986: n_2387  <= TRANSPORT a_N62_aNOT  ;
delay_1987: n_2388  <= TRANSPORT a_SCH2WRDCNTREG_F9_G  ;
and2_1988: n_2390 <=  n_2391  AND n_2392;
delay_1989: n_2391  <= TRANSPORT a_LC3_D22  ;
delay_1990: n_2392  <= TRANSPORT a_SCH2WRDCNTREG_F9_G  ;
and1_1991: n_2393 <=  gnd;
delay_1992: a_LC2_A7  <= TRANSPORT a_EQ804  ;
xor2_1993: a_EQ804 <=  n_2396  XOR n_2403;
or2_1994: n_2396 <=  n_2397  OR n_2400;
and2_1995: n_2397 <=  n_2398  AND n_2399;
delay_1996: n_2398  <= TRANSPORT a_N2560_aNOT  ;
delay_1997: n_2399  <= TRANSPORT a_LC1_A7  ;
and2_1998: n_2400 <=  n_2401  AND n_2402;
inv_1999: n_2401  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_2000: n_2402  <= TRANSPORT NOT a_LC1_A13  ;
and1_2001: n_2403 <=  gnd;
dff_2002: DFF_a8237

    PORT MAP ( D => a_EQ1058, CLK => a_SCH2WRDCNTREG_F9_G_aCLK, CLRN => a_SCH2WRDCNTREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F9_G);
inv_2003: a_SCH2WRDCNTREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2004: a_EQ1058 <=  n_2410  XOR n_2418;
or2_2005: n_2410 <=  n_2411  OR n_2414;
and2_2006: n_2411 <=  n_2412  AND n_2413;
inv_2007: n_2412  <= TRANSPORT NOT a_N2527  ;
delay_2008: n_2413  <= TRANSPORT a_LC2_A7  ;
and2_2009: n_2414 <=  n_2415  AND n_2417;
delay_2010: n_2415  <= TRANSPORT a_SCH2BWORDOUT_F9_G  ;
delay_2011: n_2417  <= TRANSPORT a_N2527  ;
and1_2012: n_2418 <=  gnd;
delay_2013: n_2419  <= TRANSPORT clk  ;
filter_2014: FILTER_a8237

    PORT MAP (IN1 => n_2419, Y => a_SCH2WRDCNTREG_F9_G_aCLK);
dff_2015: DFF_a8237

    PORT MAP ( D => a_EQ956, CLK => a_SCH1BAROUT_F9_G_aCLK, CLRN => a_SCH1BAROUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F9_G);
inv_2016: a_SCH1BAROUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2017: a_EQ956 <=  n_2428  XOR n_2435;
or2_2018: n_2428 <=  n_2429  OR n_2432;
and2_2019: n_2429 <=  n_2430  AND n_2431;
inv_2020: n_2430  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_2021: n_2431  <= TRANSPORT dbin(1)  ;
and2_2022: n_2432 <=  n_2433  AND n_2434;
delay_2023: n_2433  <= TRANSPORT a_N2585_aNOT  ;
delay_2024: n_2434  <= TRANSPORT a_SCH1BAROUT_F9_G  ;
and1_2025: n_2435 <=  gnd;
delay_2026: n_2436  <= TRANSPORT clk  ;
filter_2027: FILTER_a8237

    PORT MAP (IN1 => n_2436, Y => a_SCH1BAROUT_F9_G_aCLK);
dff_2028: DFF_a8237

    PORT MAP ( D => a_EQ1100, CLK => a_SCH3BWORDOUT_F9_G_aCLK, CLRN => a_SCH3BWORDOUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F9_G);
inv_2029: a_SCH3BWORDOUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2030: a_EQ1100 <=  n_2445  XOR n_2452;
or2_2031: n_2445 <=  n_2446  OR n_2449;
and2_2032: n_2446 <=  n_2447  AND n_2448;
inv_2033: n_2447  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_2034: n_2448  <= TRANSPORT dbin(1)  ;
and2_2035: n_2449 <=  n_2450  AND n_2451;
delay_2036: n_2450  <= TRANSPORT a_N2573_aNOT  ;
delay_2037: n_2451  <= TRANSPORT a_SCH3BWORDOUT_F9_G  ;
and1_2038: n_2452 <=  gnd;
delay_2039: n_2453  <= TRANSPORT clk  ;
filter_2040: FILTER_a8237

    PORT MAP (IN1 => n_2453, Y => a_SCH3BWORDOUT_F9_G_aCLK);
dff_2041: DFF_a8237

    PORT MAP ( D => a_EQ901, CLK => a_SCH0BWORDOUT_F2_G_aCLK, CLRN => a_SCH0BWORDOUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F2_G);
inv_2042: a_SCH0BWORDOUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2043: a_EQ901 <=  n_2462  XOR n_2469;
or2_2044: n_2462 <=  n_2463  OR n_2466;
and2_2045: n_2463 <=  n_2464  AND n_2465;
inv_2046: n_2464  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_2047: n_2465  <= TRANSPORT dbin(2)  ;
and2_2048: n_2466 <=  n_2467  AND n_2468;
delay_2049: n_2467  <= TRANSPORT a_N2578_aNOT  ;
delay_2050: n_2468  <= TRANSPORT a_SCH0BWORDOUT_F2_G  ;
and1_2051: n_2469 <=  gnd;
delay_2052: n_2470  <= TRANSPORT clk  ;
filter_2053: FILTER_a8237

    PORT MAP (IN1 => n_2470, Y => a_SCH0BWORDOUT_F2_G_aCLK);
dff_2054: DFF_a8237

    PORT MAP ( D => a_EQ1021, CLK => a_SCH2BAROUT_F10_G_aCLK, CLRN => a_SCH2BAROUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F10_G);
inv_2055: a_SCH2BAROUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2056: a_EQ1021 <=  n_2479  XOR n_2486;
or2_2057: n_2479 <=  n_2480  OR n_2483;
and2_2058: n_2480 <=  n_2481  AND n_2482;
inv_2059: n_2481  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_2060: n_2482  <= TRANSPORT dbin(2)  ;
and2_2061: n_2483 <=  n_2484  AND n_2485;
delay_2062: n_2484  <= TRANSPORT a_N2583_aNOT  ;
delay_2063: n_2485  <= TRANSPORT a_SCH2BAROUT_F10_G  ;
and1_2064: n_2486 <=  gnd;
delay_2065: n_2487  <= TRANSPORT clk  ;
filter_2066: FILTER_a8237

    PORT MAP (IN1 => n_2487, Y => a_SCH2BAROUT_F10_G_aCLK);
dff_2067: DFF_a8237

    PORT MAP ( D => a_EQ1101, CLK => a_SCH3BWORDOUT_F10_G_aCLK, CLRN => a_SCH3BWORDOUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F10_G);
inv_2068: a_SCH3BWORDOUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2069: a_EQ1101 <=  n_2496  XOR n_2503;
or2_2070: n_2496 <=  n_2497  OR n_2500;
and2_2071: n_2497 <=  n_2498  AND n_2499;
inv_2072: n_2498  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_2073: n_2499  <= TRANSPORT dbin(2)  ;
and2_2074: n_2500 <=  n_2501  AND n_2502;
delay_2075: n_2501  <= TRANSPORT a_N2573_aNOT  ;
delay_2076: n_2502  <= TRANSPORT a_SCH3BWORDOUT_F10_G  ;
and1_2077: n_2503 <=  gnd;
delay_2078: n_2504  <= TRANSPORT clk  ;
filter_2079: FILTER_a8237

    PORT MAP (IN1 => n_2504, Y => a_SCH3BWORDOUT_F10_G_aCLK);
dff_2080: DFF_a8237

    PORT MAP ( D => a_EQ1085, CLK => a_SCH3BAROUT_F10_G_aCLK, CLRN => a_SCH3BAROUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F10_G);
inv_2081: a_SCH3BAROUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2082: a_EQ1085 <=  n_2513  XOR n_2520;
or2_2083: n_2513 <=  n_2514  OR n_2517;
and2_2084: n_2514 <=  n_2515  AND n_2516;
inv_2085: n_2515  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_2086: n_2516  <= TRANSPORT dbin(2)  ;
and2_2087: n_2517 <=  n_2518  AND n_2519;
delay_2088: n_2518  <= TRANSPORT a_N2581_aNOT  ;
delay_2089: n_2519  <= TRANSPORT a_SCH3BAROUT_F10_G  ;
and1_2090: n_2520 <=  gnd;
delay_2091: n_2521  <= TRANSPORT clk  ;
filter_2092: FILTER_a8237

    PORT MAP (IN1 => n_2521, Y => a_SCH3BAROUT_F10_G_aCLK);
dff_2093: DFF_a8237

    PORT MAP ( D => a_EQ1037, CLK => a_SCH2BWORDOUT_F10_G_aCLK, CLRN => a_SCH2BWORDOUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F10_G);
inv_2094: a_SCH2BWORDOUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2095: a_EQ1037 <=  n_2530  XOR n_2541;
or3_2096: n_2530 <=  n_2531  OR n_2535  OR n_2538;
and3_2097: n_2531 <=  n_2532  AND n_2533  AND n_2534;
inv_2098: n_2532  <= TRANSPORT NOT a_LC3_D22  ;
inv_2099: n_2533  <= TRANSPORT NOT a_N62_aNOT  ;
delay_2100: n_2534  <= TRANSPORT dbin(2)  ;
and2_2101: n_2535 <=  n_2536  AND n_2537;
delay_2102: n_2536  <= TRANSPORT a_N62_aNOT  ;
delay_2103: n_2537  <= TRANSPORT a_SCH2BWORDOUT_F10_G  ;
and2_2104: n_2538 <=  n_2539  AND n_2540;
delay_2105: n_2539  <= TRANSPORT a_LC3_D22  ;
delay_2106: n_2540  <= TRANSPORT a_SCH2BWORDOUT_F10_G  ;
and1_2107: n_2541 <=  gnd;
delay_2108: n_2542  <= TRANSPORT clk  ;
filter_2109: FILTER_a8237

    PORT MAP (IN1 => n_2542, Y => a_SCH2BWORDOUT_F10_G_aCLK);
dff_2110: DFF_a8237

    PORT MAP ( D => a_EQ957, CLK => a_SCH1BAROUT_F10_G_aCLK, CLRN => a_SCH1BAROUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F10_G);
inv_2111: a_SCH1BAROUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2112: a_EQ957 <=  n_2551  XOR n_2558;
or2_2113: n_2551 <=  n_2552  OR n_2555;
and2_2114: n_2552 <=  n_2553  AND n_2554;
inv_2115: n_2553  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_2116: n_2554  <= TRANSPORT dbin(2)  ;
and2_2117: n_2555 <=  n_2556  AND n_2557;
delay_2118: n_2556  <= TRANSPORT a_N2585_aNOT  ;
delay_2119: n_2557  <= TRANSPORT a_SCH1BAROUT_F10_G  ;
and1_2120: n_2558 <=  gnd;
delay_2121: n_2559  <= TRANSPORT clk  ;
filter_2122: FILTER_a8237

    PORT MAP (IN1 => n_2559, Y => a_SCH1BAROUT_F10_G_aCLK);
dff_2123: DFF_a8237

    PORT MAP ( D => a_EQ909, CLK => a_SCH0BWORDOUT_F10_G_aCLK, CLRN => a_SCH0BWORDOUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F10_G);
inv_2124: a_SCH0BWORDOUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2125: a_EQ909 <=  n_2568  XOR n_2579;
or3_2126: n_2568 <=  n_2569  OR n_2573  OR n_2576;
and3_2127: n_2569 <=  n_2570  AND n_2571  AND n_2572;
inv_2128: n_2570  <= TRANSPORT NOT a_LC3_D22  ;
inv_2129: n_2571  <= TRANSPORT NOT a_N2353  ;
delay_2130: n_2572  <= TRANSPORT dbin(2)  ;
and2_2131: n_2573 <=  n_2574  AND n_2575;
delay_2132: n_2574  <= TRANSPORT a_N2353  ;
delay_2133: n_2575  <= TRANSPORT a_SCH0BWORDOUT_F10_G  ;
and2_2134: n_2576 <=  n_2577  AND n_2578;
delay_2135: n_2577  <= TRANSPORT a_LC3_D22  ;
delay_2136: n_2578  <= TRANSPORT a_SCH0BWORDOUT_F10_G  ;
and1_2137: n_2579 <=  gnd;
delay_2138: n_2580  <= TRANSPORT clk  ;
filter_2139: FILTER_a8237

    PORT MAP (IN1 => n_2580, Y => a_SCH0BWORDOUT_F10_G_aCLK);
dff_2140: DFF_a8237

    PORT MAP ( D => a_EQ893, CLK => a_SCH0BAROUT_F10_G_aCLK, CLRN => a_SCH0BAROUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F10_G);
inv_2141: a_SCH0BAROUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2142: a_EQ893 <=  n_2589  XOR n_2596;
or2_2143: n_2589 <=  n_2590  OR n_2593;
and2_2144: n_2590 <=  n_2591  AND n_2592;
delay_2145: n_2591  <= TRANSPORT a_N2587_aNOT  ;
delay_2146: n_2592  <= TRANSPORT a_SCH0BAROUT_F10_G  ;
and2_2147: n_2593 <=  n_2594  AND n_2595;
inv_2148: n_2594  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_2149: n_2595  <= TRANSPORT dbin(2)  ;
and1_2150: n_2596 <=  gnd;
delay_2151: n_2597  <= TRANSPORT clk  ;
filter_2152: FILTER_a8237

    PORT MAP (IN1 => n_2597, Y => a_SCH0BAROUT_F10_G_aCLK);
dff_2153: DFF_a8237

    PORT MAP ( D => a_EQ1022, CLK => a_SCH2BAROUT_F11_G_aCLK, CLRN => a_SCH2BAROUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F11_G);
inv_2154: a_SCH2BAROUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2155: a_EQ1022 <=  n_2606  XOR n_2613;
or2_2156: n_2606 <=  n_2607  OR n_2610;
and2_2157: n_2607 <=  n_2608  AND n_2609;
inv_2158: n_2608  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_2159: n_2609  <= TRANSPORT dbin(3)  ;
and2_2160: n_2610 <=  n_2611  AND n_2612;
delay_2161: n_2611  <= TRANSPORT a_N2583_aNOT  ;
delay_2162: n_2612  <= TRANSPORT a_SCH2BAROUT_F11_G  ;
and1_2163: n_2613 <=  gnd;
delay_2164: n_2614  <= TRANSPORT clk  ;
filter_2165: FILTER_a8237

    PORT MAP (IN1 => n_2614, Y => a_SCH2BAROUT_F11_G_aCLK);
dff_2166: DFF_a8237

    PORT MAP ( D => a_EQ1086, CLK => a_SCH3BAROUT_F11_G_aCLK, CLRN => a_SCH3BAROUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F11_G);
inv_2167: a_SCH3BAROUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2168: a_EQ1086 <=  n_2623  XOR n_2630;
or2_2169: n_2623 <=  n_2624  OR n_2627;
and2_2170: n_2624 <=  n_2625  AND n_2626;
inv_2171: n_2625  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_2172: n_2626  <= TRANSPORT dbin(3)  ;
and2_2173: n_2627 <=  n_2628  AND n_2629;
delay_2174: n_2628  <= TRANSPORT a_N2581_aNOT  ;
delay_2175: n_2629  <= TRANSPORT a_SCH3BAROUT_F11_G  ;
and1_2176: n_2630 <=  gnd;
delay_2177: n_2631  <= TRANSPORT clk  ;
filter_2178: FILTER_a8237

    PORT MAP (IN1 => n_2631, Y => a_SCH3BAROUT_F11_G_aCLK);
dff_2179: DFF_a8237

    PORT MAP ( D => a_EQ894, CLK => a_SCH0BAROUT_F11_G_aCLK, CLRN => a_SCH0BAROUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F11_G);
inv_2180: a_SCH0BAROUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2181: a_EQ894 <=  n_2640  XOR n_2647;
or2_2182: n_2640 <=  n_2641  OR n_2644;
and2_2183: n_2641 <=  n_2642  AND n_2643;
inv_2184: n_2642  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_2185: n_2643  <= TRANSPORT dbin(3)  ;
and2_2186: n_2644 <=  n_2645  AND n_2646;
delay_2187: n_2645  <= TRANSPORT a_N2587_aNOT  ;
delay_2188: n_2646  <= TRANSPORT a_SCH0BAROUT_F11_G  ;
and1_2189: n_2647 <=  gnd;
delay_2190: n_2648  <= TRANSPORT clk  ;
filter_2191: FILTER_a8237

    PORT MAP (IN1 => n_2648, Y => a_SCH0BAROUT_F11_G_aCLK);
dff_2192: DFF_a8237

    PORT MAP ( D => a_EQ958, CLK => a_SCH1BAROUT_F11_G_aCLK, CLRN => a_SCH1BAROUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F11_G);
inv_2193: a_SCH1BAROUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2194: a_EQ958 <=  n_2657  XOR n_2664;
or2_2195: n_2657 <=  n_2658  OR n_2661;
and2_2196: n_2658 <=  n_2659  AND n_2660;
inv_2197: n_2659  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_2198: n_2660  <= TRANSPORT dbin(3)  ;
and2_2199: n_2661 <=  n_2662  AND n_2663;
delay_2200: n_2662  <= TRANSPORT a_N2585_aNOT  ;
delay_2201: n_2663  <= TRANSPORT a_SCH1BAROUT_F11_G  ;
and1_2202: n_2664 <=  gnd;
delay_2203: n_2665  <= TRANSPORT clk  ;
filter_2204: FILTER_a8237

    PORT MAP (IN1 => n_2665, Y => a_SCH1BAROUT_F11_G_aCLK);
delay_2205: a_LC1_C10  <= TRANSPORT a_EQ767  ;
xor2_2206: a_EQ767 <=  n_2669  XOR n_2676;
or2_2207: n_2669 <=  n_2670  OR n_2673;
and2_2208: n_2670 <=  n_2671  AND n_2672;
inv_2209: n_2671  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_2210: n_2672  <= TRANSPORT dbin(3)  ;
and2_2211: n_2673 <=  n_2674  AND n_2675;
delay_2212: n_2674  <= TRANSPORT a_N2578_aNOT  ;
delay_2213: n_2675  <= TRANSPORT a_SCH0WRDCNTREG_F3_G  ;
and1_2214: n_2676 <=  gnd;
delay_2215: a_LC3_C10  <= TRANSPORT a_EQ768  ;
xor2_2216: a_EQ768 <=  n_2679  XOR n_2686;
or2_2217: n_2679 <=  n_2680  OR n_2683;
and2_2218: n_2680 <=  n_2681  AND n_2682;
inv_2219: n_2681  <= TRANSPORT NOT a_LC1_C21  ;
inv_2220: n_2682  <= TRANSPORT NOT a_N2558_aNOT  ;
and2_2221: n_2683 <=  n_2684  AND n_2685;
delay_2222: n_2684  <= TRANSPORT a_N2558_aNOT  ;
delay_2223: n_2685  <= TRANSPORT a_LC1_C10  ;
and1_2224: n_2686 <=  gnd;
dff_2225: DFF_a8237

    PORT MAP ( D => a_EQ924, CLK => a_SCH0WRDCNTREG_F3_G_aCLK, CLRN => a_SCH0WRDCNTREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F3_G);
inv_2226: a_SCH0WRDCNTREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2227: a_EQ924 <=  n_2693  XOR n_2701;
or2_2228: n_2693 <=  n_2694  OR n_2697;
and2_2229: n_2694 <=  n_2695  AND n_2696;
inv_2230: n_2695  <= TRANSPORT NOT a_N2525  ;
delay_2231: n_2696  <= TRANSPORT a_LC3_C10  ;
and2_2232: n_2697 <=  n_2698  AND n_2700;
delay_2233: n_2698  <= TRANSPORT a_SCH0BWORDOUT_F3_G  ;
delay_2234: n_2700  <= TRANSPORT a_N2525  ;
and1_2235: n_2701 <=  gnd;
delay_2236: n_2702  <= TRANSPORT clk  ;
filter_2237: FILTER_a8237

    PORT MAP (IN1 => n_2702, Y => a_SCH0WRDCNTREG_F3_G_aCLK);
delay_2238: a_LC2_C22  <= TRANSPORT a_EQ790  ;
xor2_2239: a_EQ790 <=  n_2706  XOR n_2713;
or2_2240: n_2706 <=  n_2707  OR n_2710;
and2_2241: n_2707 <=  n_2708  AND n_2709;
inv_2242: n_2708  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_2243: n_2709  <= TRANSPORT dbin(3)  ;
and2_2244: n_2710 <=  n_2711  AND n_2712;
delay_2245: n_2711  <= TRANSPORT a_N2576_aNOT  ;
delay_2246: n_2712  <= TRANSPORT a_SCH1WRDCNTREG_F3_G  ;
and1_2247: n_2713 <=  gnd;
delay_2248: a_LC5_C22  <= TRANSPORT a_EQ791  ;
xor2_2249: a_EQ791 <=  n_2716  XOR n_2723;
or2_2250: n_2716 <=  n_2717  OR n_2720;
and2_2251: n_2717 <=  n_2718  AND n_2719;
inv_2252: n_2718  <= TRANSPORT NOT a_LC1_C21  ;
inv_2253: n_2719  <= TRANSPORT NOT a_N2559_aNOT  ;
and2_2254: n_2720 <=  n_2721  AND n_2722;
delay_2255: n_2721  <= TRANSPORT a_N2559_aNOT  ;
delay_2256: n_2722  <= TRANSPORT a_LC2_C22  ;
and1_2257: n_2723 <=  gnd;
dff_2258: DFF_a8237

    PORT MAP ( D => a_EQ988, CLK => a_SCH1WRDCNTREG_F3_G_aCLK, CLRN => a_SCH1WRDCNTREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F3_G);
inv_2259: a_SCH1WRDCNTREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2260: a_EQ988 <=  n_2730  XOR n_2738;
or2_2261: n_2730 <=  n_2731  OR n_2734;
and2_2262: n_2731 <=  n_2732  AND n_2733;
inv_2263: n_2732  <= TRANSPORT NOT a_N2526  ;
delay_2264: n_2733  <= TRANSPORT a_LC5_C22  ;
and2_2265: n_2734 <=  n_2735  AND n_2737;
delay_2266: n_2735  <= TRANSPORT a_SCH1BWORDOUT_F3_G  ;
delay_2267: n_2737  <= TRANSPORT a_N2526  ;
and1_2268: n_2738 <=  gnd;
delay_2269: n_2739  <= TRANSPORT clk  ;
filter_2270: FILTER_a8237

    PORT MAP (IN1 => n_2739, Y => a_SCH1WRDCNTREG_F3_G_aCLK);
delay_2271: a_LC2_C7  <= TRANSPORT a_EQ810  ;
xor2_2272: a_EQ810 <=  n_2743  XOR n_2752;
or2_2273: n_2743 <=  n_2744  OR n_2748;
and3_2274: n_2744 <=  n_2745  AND n_2746  AND n_2747;
inv_2275: n_2745  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_2276: n_2746  <= TRANSPORT a_N756  ;
delay_2277: n_2747  <= TRANSPORT dbin(3)  ;
and3_2278: n_2748 <=  n_2749  AND n_2750  AND n_2751;
delay_2279: n_2749  <= TRANSPORT a_N2574_aNOT  ;
delay_2280: n_2750  <= TRANSPORT a_N756  ;
delay_2281: n_2751  <= TRANSPORT a_SCH2WRDCNTREG_F3_G  ;
and1_2282: n_2752 <=  gnd;
delay_2283: a_N808  <= TRANSPORT a_N808_aIN  ;
xor2_2284: a_N808_aIN <=  n_2755  XOR n_2759;
or1_2285: n_2755 <=  n_2756;
and2_2286: n_2756 <=  n_2757  AND n_2758;
inv_2287: n_2757  <= TRANSPORT NOT a_LC1_C21  ;
delay_2288: n_2758  <= TRANSPORT a_N858  ;
and1_2289: n_2759 <=  gnd;
dff_2290: DFF_a8237

    PORT MAP ( D => a_EQ1052, CLK => a_SCH2WRDCNTREG_F3_G_aCLK, CLRN => a_SCH2WRDCNTREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F3_G);
inv_2291: a_SCH2WRDCNTREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2292: a_EQ1052 <=  n_2766  XOR n_2774;
or3_2293: n_2766 <=  n_2767  OR n_2769  OR n_2771;
and1_2294: n_2767 <=  n_2768;
delay_2295: n_2768  <= TRANSPORT a_LC2_C7  ;
and1_2296: n_2769 <=  n_2770;
delay_2297: n_2770  <= TRANSPORT a_N808  ;
and2_2298: n_2771 <=  n_2772  AND n_2773;
delay_2299: n_2772  <= TRANSPORT a_SCH2BWORDOUT_F3_G  ;
delay_2300: n_2773  <= TRANSPORT a_N2527  ;
and1_2301: n_2774 <=  gnd;
delay_2302: n_2775  <= TRANSPORT clk  ;
filter_2303: FILTER_a8237

    PORT MAP (IN1 => n_2775, Y => a_SCH2WRDCNTREG_F3_G_aCLK);
dff_2304: DFF_a8237

    PORT MAP ( D => a_EQ1094, CLK => a_SCH3BWORDOUT_F3_G_aCLK, CLRN => a_SCH3BWORDOUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F3_G);
inv_2305: a_SCH3BWORDOUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2306: a_EQ1094 <=  n_2784  XOR n_2791;
or2_2307: n_2784 <=  n_2785  OR n_2788;
and2_2308: n_2785 <=  n_2786  AND n_2787;
inv_2309: n_2786  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_2310: n_2787  <= TRANSPORT dbin(3)  ;
and2_2311: n_2788 <=  n_2789  AND n_2790;
delay_2312: n_2789  <= TRANSPORT a_N2572_aNOT  ;
delay_2313: n_2790  <= TRANSPORT a_SCH3BWORDOUT_F3_G  ;
and1_2314: n_2791 <=  gnd;
delay_2315: n_2792  <= TRANSPORT clk  ;
filter_2316: FILTER_a8237

    PORT MAP (IN1 => n_2792, Y => a_SCH3BWORDOUT_F3_G_aCLK);
delay_2317: a_LC1_C3  <= TRANSPORT a_EQ765  ;
xor2_2318: a_EQ765 <=  n_2796  XOR n_2804;
or2_2319: n_2796 <=  n_2797  OR n_2800;
and2_2320: n_2797 <=  n_2798  AND n_2799;
inv_2321: n_2798  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_2322: n_2799  <= TRANSPORT dbin(4)  ;
and2_2323: n_2800 <=  n_2801  AND n_2802;
delay_2324: n_2801  <= TRANSPORT a_N2578_aNOT  ;
delay_2325: n_2802  <= TRANSPORT a_SCH0WRDCNTREG_F4_G  ;
and1_2326: n_2804 <=  gnd;
delay_2327: a_LC2_C3  <= TRANSPORT a_EQ766  ;
xor2_2328: a_EQ766 <=  n_2807  XOR n_2819;
or3_2329: n_2807 <=  n_2808  OR n_2811  OR n_2815;
and2_2330: n_2808 <=  n_2809  AND n_2810;
delay_2331: n_2809  <= TRANSPORT a_N2558_aNOT  ;
delay_2332: n_2810  <= TRANSPORT a_LC1_C3  ;
and3_2333: n_2811 <=  n_2812  AND n_2813  AND n_2814;
delay_2334: n_2812  <= TRANSPORT a_LC3_C13  ;
inv_2335: n_2813  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_2336: n_2814  <= TRANSPORT a_N3552  ;
and3_2337: n_2815 <=  n_2816  AND n_2817  AND n_2818;
inv_2338: n_2816  <= TRANSPORT NOT a_LC3_C13  ;
inv_2339: n_2817  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_2340: n_2818  <= TRANSPORT NOT a_N3552  ;
and1_2341: n_2819 <=  gnd;
dff_2342: DFF_a8237

    PORT MAP ( D => a_EQ925, CLK => a_SCH0WRDCNTREG_F4_G_aCLK, CLRN => a_SCH0WRDCNTREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F4_G);
inv_2343: a_SCH0WRDCNTREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2344: a_EQ925 <=  n_2826  XOR n_2833;
or2_2345: n_2826 <=  n_2827  OR n_2830;
and2_2346: n_2827 <=  n_2828  AND n_2829;
inv_2347: n_2828  <= TRANSPORT NOT a_N2525  ;
delay_2348: n_2829  <= TRANSPORT a_LC2_C3  ;
and2_2349: n_2830 <=  n_2831  AND n_2832;
delay_2350: n_2831  <= TRANSPORT a_SCH0BWORDOUT_F4_G  ;
delay_2351: n_2832  <= TRANSPORT a_N2525  ;
and1_2352: n_2833 <=  gnd;
delay_2353: n_2834  <= TRANSPORT clk  ;
filter_2354: FILTER_a8237

    PORT MAP (IN1 => n_2834, Y => a_SCH0WRDCNTREG_F4_G_aCLK);
delay_2355: a_LC2_C1  <= TRANSPORT a_EQ829  ;
xor2_2356: a_EQ829 <=  n_2838  XOR n_2848;
or2_2357: n_2838 <=  n_2839  OR n_2843;
and3_2358: n_2839 <=  n_2840  AND n_2841  AND n_2842;
inv_2359: n_2840  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_2360: n_2841  <= TRANSPORT a_N1095  ;
delay_2361: n_2842  <= TRANSPORT dbin(4)  ;
and3_2362: n_2843 <=  n_2844  AND n_2845  AND n_2846;
delay_2363: n_2844  <= TRANSPORT a_N2572_aNOT  ;
delay_2364: n_2845  <= TRANSPORT a_N1095  ;
delay_2365: n_2846  <= TRANSPORT a_SCH3WRDCNTREG_F4_G  ;
and1_2366: n_2848 <=  gnd;
delay_2367: a_N1037_aNOT  <= TRANSPORT a_EQ344  ;
xor2_2368: a_EQ344 <=  n_2851  XOR n_2860;
or2_2369: n_2851 <=  n_2852  OR n_2856;
and3_2370: n_2852 <=  n_2853  AND n_2854  AND n_2855;
delay_2371: n_2853  <= TRANSPORT a_LC3_C13  ;
delay_2372: n_2854  <= TRANSPORT a_N1094  ;
delay_2373: n_2855  <= TRANSPORT a_N3552  ;
and3_2374: n_2856 <=  n_2857  AND n_2858  AND n_2859;
inv_2375: n_2857  <= TRANSPORT NOT a_LC3_C13  ;
delay_2376: n_2858  <= TRANSPORT a_N1094  ;
inv_2377: n_2859  <= TRANSPORT NOT a_N3552  ;
and1_2378: n_2860 <=  gnd;
dff_2379: DFF_a8237

    PORT MAP ( D => a_EQ1117, CLK => a_SCH3WRDCNTREG_F4_G_aCLK, CLRN => a_SCH3WRDCNTREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F4_G);
inv_2380: a_SCH3WRDCNTREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2381: a_EQ1117 <=  n_2867  XOR n_2875;
or3_2382: n_2867 <=  n_2868  OR n_2870  OR n_2872;
and1_2383: n_2868 <=  n_2869;
delay_2384: n_2869  <= TRANSPORT a_LC2_C1  ;
and1_2385: n_2870 <=  n_2871;
delay_2386: n_2871  <= TRANSPORT a_N1037_aNOT  ;
and2_2387: n_2872 <=  n_2873  AND n_2874;
delay_2388: n_2873  <= TRANSPORT a_SCH3BWORDOUT_F4_G  ;
delay_2389: n_2874  <= TRANSPORT a_N2528  ;
and1_2390: n_2875 <=  gnd;
delay_2391: n_2876  <= TRANSPORT clk  ;
filter_2392: FILTER_a8237

    PORT MAP (IN1 => n_2876, Y => a_SCH3WRDCNTREG_F4_G_aCLK);
delay_2393: a_LC4_C18  <= TRANSPORT a_EQ809  ;
xor2_2394: a_EQ809 <=  n_2880  XOR n_2890;
or2_2395: n_2880 <=  n_2881  OR n_2885;
and3_2396: n_2881 <=  n_2882  AND n_2883  AND n_2884;
inv_2397: n_2882  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_2398: n_2883  <= TRANSPORT a_N756  ;
delay_2399: n_2884  <= TRANSPORT dbin(4)  ;
and3_2400: n_2885 <=  n_2886  AND n_2887  AND n_2888;
delay_2401: n_2886  <= TRANSPORT a_N2574_aNOT  ;
delay_2402: n_2887  <= TRANSPORT a_N756  ;
delay_2403: n_2888  <= TRANSPORT a_SCH2WRDCNTREG_F4_G  ;
and1_2404: n_2890 <=  gnd;
delay_2405: a_N815  <= TRANSPORT a_EQ304  ;
xor2_2406: a_EQ304 <=  n_2893  XOR n_2902;
or2_2407: n_2893 <=  n_2894  OR n_2898;
and3_2408: n_2894 <=  n_2895  AND n_2896  AND n_2897;
delay_2409: n_2895  <= TRANSPORT a_LC3_C13  ;
delay_2410: n_2896  <= TRANSPORT a_N858  ;
delay_2411: n_2897  <= TRANSPORT a_N3552  ;
and3_2412: n_2898 <=  n_2899  AND n_2900  AND n_2901;
inv_2413: n_2899  <= TRANSPORT NOT a_LC3_C13  ;
delay_2414: n_2900  <= TRANSPORT a_N858  ;
inv_2415: n_2901  <= TRANSPORT NOT a_N3552  ;
and1_2416: n_2902 <=  gnd;
dff_2417: DFF_a8237

    PORT MAP ( D => a_EQ1053, CLK => a_SCH2WRDCNTREG_F4_G_aCLK, CLRN => a_SCH2WRDCNTREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F4_G);
inv_2418: a_SCH2WRDCNTREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2419: a_EQ1053 <=  n_2909  XOR n_2917;
or3_2420: n_2909 <=  n_2910  OR n_2912  OR n_2914;
and1_2421: n_2910 <=  n_2911;
delay_2422: n_2911  <= TRANSPORT a_LC4_C18  ;
and1_2423: n_2912 <=  n_2913;
delay_2424: n_2913  <= TRANSPORT a_N815  ;
and2_2425: n_2914 <=  n_2915  AND n_2916;
delay_2426: n_2915  <= TRANSPORT a_SCH2BWORDOUT_F4_G  ;
delay_2427: n_2916  <= TRANSPORT a_N2527  ;
and1_2428: n_2917 <=  gnd;
delay_2429: n_2918  <= TRANSPORT clk  ;
filter_2430: FILTER_a8237

    PORT MAP (IN1 => n_2918, Y => a_SCH2WRDCNTREG_F4_G_aCLK);
delay_2431: a_LC5_F4  <= TRANSPORT a_EQ788  ;
xor2_2432: a_EQ788 <=  n_2922  XOR n_2930;
or2_2433: n_2922 <=  n_2923  OR n_2926;
and2_2434: n_2923 <=  n_2924  AND n_2925;
inv_2435: n_2924  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_2436: n_2925  <= TRANSPORT dbin(4)  ;
and2_2437: n_2926 <=  n_2927  AND n_2928;
delay_2438: n_2927  <= TRANSPORT a_N2576_aNOT  ;
delay_2439: n_2928  <= TRANSPORT a_SCH1WRDCNTREG_F4_G  ;
and1_2440: n_2930 <=  gnd;
delay_2441: a_LC6_F4  <= TRANSPORT a_EQ789  ;
xor2_2442: a_EQ789 <=  n_2933  XOR n_2945;
or3_2443: n_2933 <=  n_2934  OR n_2937  OR n_2941;
and2_2444: n_2934 <=  n_2935  AND n_2936;
delay_2445: n_2935  <= TRANSPORT a_N2559_aNOT  ;
delay_2446: n_2936  <= TRANSPORT a_LC5_F4  ;
and3_2447: n_2937 <=  n_2938  AND n_2939  AND n_2940;
delay_2448: n_2938  <= TRANSPORT a_LC3_C13  ;
inv_2449: n_2939  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_2450: n_2940  <= TRANSPORT a_N3552  ;
and3_2451: n_2941 <=  n_2942  AND n_2943  AND n_2944;
inv_2452: n_2942  <= TRANSPORT NOT a_LC3_C13  ;
inv_2453: n_2943  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_2454: n_2944  <= TRANSPORT NOT a_N3552  ;
and1_2455: n_2945 <=  gnd;
dff_2456: DFF_a8237

    PORT MAP ( D => a_EQ989, CLK => a_SCH1WRDCNTREG_F4_G_aCLK, CLRN => a_SCH1WRDCNTREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F4_G);
inv_2457: a_SCH1WRDCNTREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2458: a_EQ989 <=  n_2952  XOR n_2959;
or2_2459: n_2952 <=  n_2953  OR n_2956;
and2_2460: n_2953 <=  n_2954  AND n_2955;
inv_2461: n_2954  <= TRANSPORT NOT a_N2526  ;
delay_2462: n_2955  <= TRANSPORT a_LC6_F4  ;
and2_2463: n_2956 <=  n_2957  AND n_2958;
delay_2464: n_2957  <= TRANSPORT a_SCH1BWORDOUT_F4_G  ;
delay_2465: n_2958  <= TRANSPORT a_N2526  ;
and1_2466: n_2959 <=  gnd;
delay_2467: n_2960  <= TRANSPORT clk  ;
filter_2468: FILTER_a8237

    PORT MAP (IN1 => n_2960, Y => a_SCH1WRDCNTREG_F4_G_aCLK);
dff_2469: DFF_a8237

    PORT MAP ( D => a_EQ1023, CLK => a_SCH2BAROUT_F12_G_aCLK, CLRN => a_SCH2BAROUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F12_G);
inv_2470: a_SCH2BAROUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2471: a_EQ1023 <=  n_2969  XOR n_2976;
or2_2472: n_2969 <=  n_2970  OR n_2973;
and2_2473: n_2970 <=  n_2971  AND n_2972;
inv_2474: n_2971  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_2475: n_2972  <= TRANSPORT dbin(4)  ;
and2_2476: n_2973 <=  n_2974  AND n_2975;
delay_2477: n_2974  <= TRANSPORT a_N2583_aNOT  ;
delay_2478: n_2975  <= TRANSPORT a_SCH2BAROUT_F12_G  ;
and1_2479: n_2976 <=  gnd;
delay_2480: n_2977  <= TRANSPORT clk  ;
filter_2481: FILTER_a8237

    PORT MAP (IN1 => n_2977, Y => a_SCH2BAROUT_F12_G_aCLK);
dff_2482: DFF_a8237

    PORT MAP ( D => a_EQ895, CLK => a_SCH0BAROUT_F12_G_aCLK, CLRN => a_SCH0BAROUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F12_G);
inv_2483: a_SCH0BAROUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2484: a_EQ895 <=  n_2986  XOR n_2993;
or2_2485: n_2986 <=  n_2987  OR n_2990;
and2_2486: n_2987 <=  n_2988  AND n_2989;
inv_2487: n_2988  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_2488: n_2989  <= TRANSPORT dbin(4)  ;
and2_2489: n_2990 <=  n_2991  AND n_2992;
delay_2490: n_2991  <= TRANSPORT a_N2587_aNOT  ;
delay_2491: n_2992  <= TRANSPORT a_SCH0BAROUT_F12_G  ;
and1_2492: n_2993 <=  gnd;
delay_2493: n_2994  <= TRANSPORT clk  ;
filter_2494: FILTER_a8237

    PORT MAP (IN1 => n_2994, Y => a_SCH0BAROUT_F12_G_aCLK);
dff_2495: DFF_a8237

    PORT MAP ( D => a_EQ1087, CLK => a_SCH3BAROUT_F12_G_aCLK, CLRN => a_SCH3BAROUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F12_G);
inv_2496: a_SCH3BAROUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2497: a_EQ1087 <=  n_3003  XOR n_3010;
or2_2498: n_3003 <=  n_3004  OR n_3007;
and2_2499: n_3004 <=  n_3005  AND n_3006;
inv_2500: n_3005  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_2501: n_3006  <= TRANSPORT dbin(4)  ;
and2_2502: n_3007 <=  n_3008  AND n_3009;
delay_2503: n_3008  <= TRANSPORT a_N2581_aNOT  ;
delay_2504: n_3009  <= TRANSPORT a_SCH3BAROUT_F12_G  ;
and1_2505: n_3010 <=  gnd;
delay_2506: n_3011  <= TRANSPORT clk  ;
filter_2507: FILTER_a8237

    PORT MAP (IN1 => n_3011, Y => a_SCH3BAROUT_F12_G_aCLK);
dff_2508: DFF_a8237

    PORT MAP ( D => a_EQ904, CLK => a_SCH0BWORDOUT_F5_G_aCLK, CLRN => a_SCH0BWORDOUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F5_G);
inv_2509: a_SCH0BWORDOUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2510: a_EQ904 <=  n_3020  XOR n_3027;
or2_2511: n_3020 <=  n_3021  OR n_3024;
and2_2512: n_3021 <=  n_3022  AND n_3023;
inv_2513: n_3022  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_2514: n_3023  <= TRANSPORT dbin(5)  ;
and2_2515: n_3024 <=  n_3025  AND n_3026;
delay_2516: n_3025  <= TRANSPORT a_N2578_aNOT  ;
delay_2517: n_3026  <= TRANSPORT a_SCH0BWORDOUT_F5_G  ;
and1_2518: n_3027 <=  gnd;
delay_2519: n_3028  <= TRANSPORT clk  ;
filter_2520: FILTER_a8237

    PORT MAP (IN1 => n_3028, Y => a_SCH0BWORDOUT_F5_G_aCLK);
dff_2521: DFF_a8237

    PORT MAP ( D => a_EQ1096, CLK => a_SCH3BWORDOUT_F5_G_aCLK, CLRN => a_SCH3BWORDOUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F5_G);
inv_2522: a_SCH3BWORDOUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2523: a_EQ1096 <=  n_3037  XOR n_3044;
or2_2524: n_3037 <=  n_3038  OR n_3041;
and2_2525: n_3038 <=  n_3039  AND n_3040;
inv_2526: n_3039  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_2527: n_3040  <= TRANSPORT dbin(5)  ;
and2_2528: n_3041 <=  n_3042  AND n_3043;
delay_2529: n_3042  <= TRANSPORT a_N2572_aNOT  ;
delay_2530: n_3043  <= TRANSPORT a_SCH3BWORDOUT_F5_G  ;
and1_2531: n_3044 <=  gnd;
delay_2532: n_3045  <= TRANSPORT clk  ;
filter_2533: FILTER_a8237

    PORT MAP (IN1 => n_3045, Y => a_SCH3BWORDOUT_F5_G_aCLK);
dff_2534: DFF_a8237

    PORT MAP ( D => a_EQ968, CLK => a_SCH1BWORDOUT_F5_G_aCLK, CLRN => a_SCH1BWORDOUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F5_G);
inv_2535: a_SCH1BWORDOUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2536: a_EQ968 <=  n_3054  XOR n_3061;
or2_2537: n_3054 <=  n_3055  OR n_3058;
and2_2538: n_3055 <=  n_3056  AND n_3057;
inv_2539: n_3056  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_2540: n_3057  <= TRANSPORT dbin(5)  ;
and2_2541: n_3058 <=  n_3059  AND n_3060;
delay_2542: n_3059  <= TRANSPORT a_N2576_aNOT  ;
delay_2543: n_3060  <= TRANSPORT a_SCH1BWORDOUT_F5_G  ;
and1_2544: n_3061 <=  gnd;
delay_2545: n_3062  <= TRANSPORT clk  ;
filter_2546: FILTER_a8237

    PORT MAP (IN1 => n_3062, Y => a_SCH1BWORDOUT_F5_G_aCLK);
dff_2547: DFF_a8237

    PORT MAP ( D => a_EQ1032, CLK => a_SCH2BWORDOUT_F5_G_aCLK, CLRN => a_SCH2BWORDOUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F5_G);
inv_2548: a_SCH2BWORDOUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2549: a_EQ1032 <=  n_3071  XOR n_3078;
or2_2550: n_3071 <=  n_3072  OR n_3075;
and2_2551: n_3072 <=  n_3073  AND n_3074;
inv_2552: n_3073  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_2553: n_3074  <= TRANSPORT dbin(5)  ;
and2_2554: n_3075 <=  n_3076  AND n_3077;
delay_2555: n_3076  <= TRANSPORT a_N2574_aNOT  ;
delay_2556: n_3077  <= TRANSPORT a_SCH2BWORDOUT_F5_G  ;
and1_2557: n_3078 <=  gnd;
delay_2558: n_3079  <= TRANSPORT clk  ;
filter_2559: FILTER_a8237

    PORT MAP (IN1 => n_3079, Y => a_SCH2BWORDOUT_F5_G_aCLK);
dff_2560: DFF_a8237

    PORT MAP ( D => a_EQ912, CLK => a_SCH0BWORDOUT_F13_G_aCLK, CLRN => a_SCH0BWORDOUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F13_G);
inv_2561: a_SCH0BWORDOUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2562: a_EQ912 <=  n_3088  XOR n_3099;
or3_2563: n_3088 <=  n_3089  OR n_3093  OR n_3096;
and3_2564: n_3089 <=  n_3090  AND n_3091  AND n_3092;
inv_2565: n_3090  <= TRANSPORT NOT a_LC3_D22  ;
inv_2566: n_3091  <= TRANSPORT NOT a_N2353  ;
delay_2567: n_3092  <= TRANSPORT dbin(5)  ;
and2_2568: n_3093 <=  n_3094  AND n_3095;
delay_2569: n_3094  <= TRANSPORT a_N2353  ;
delay_2570: n_3095  <= TRANSPORT a_SCH0BWORDOUT_F13_G  ;
and2_2571: n_3096 <=  n_3097  AND n_3098;
delay_2572: n_3097  <= TRANSPORT a_LC3_D22  ;
delay_2573: n_3098  <= TRANSPORT a_SCH0BWORDOUT_F13_G  ;
and1_2574: n_3099 <=  gnd;
delay_2575: n_3100  <= TRANSPORT clk  ;
filter_2576: FILTER_a8237

    PORT MAP (IN1 => n_3100, Y => a_SCH0BWORDOUT_F13_G_aCLK);
dff_2577: DFF_a8237

    PORT MAP ( D => a_EQ1104, CLK => a_SCH3BWORDOUT_F13_G_aCLK, CLRN => a_SCH3BWORDOUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F13_G);
inv_2578: a_SCH3BWORDOUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2579: a_EQ1104 <=  n_3109  XOR n_3116;
or2_2580: n_3109 <=  n_3110  OR n_3113;
and2_2581: n_3110 <=  n_3111  AND n_3112;
inv_2582: n_3111  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_2583: n_3112  <= TRANSPORT dbin(5)  ;
and2_2584: n_3113 <=  n_3114  AND n_3115;
delay_2585: n_3114  <= TRANSPORT a_N2573_aNOT  ;
delay_2586: n_3115  <= TRANSPORT a_SCH3BWORDOUT_F13_G  ;
and1_2587: n_3116 <=  gnd;
delay_2588: n_3117  <= TRANSPORT clk  ;
filter_2589: FILTER_a8237

    PORT MAP (IN1 => n_3117, Y => a_SCH3BWORDOUT_F13_G_aCLK);
dff_2590: DFF_a8237

    PORT MAP ( D => a_EQ976, CLK => a_SCH1BWORDOUT_F13_G_aCLK, CLRN => a_SCH1BWORDOUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F13_G);
inv_2591: a_SCH1BWORDOUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2592: a_EQ976 <=  n_3126  XOR n_3133;
or2_2593: n_3126 <=  n_3127  OR n_3130;
and2_2594: n_3127 <=  n_3128  AND n_3129;
inv_2595: n_3128  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_2596: n_3129  <= TRANSPORT dbin(5)  ;
and2_2597: n_3130 <=  n_3131  AND n_3132;
delay_2598: n_3131  <= TRANSPORT a_N2577_aNOT  ;
delay_2599: n_3132  <= TRANSPORT a_SCH1BWORDOUT_F13_G  ;
and1_2600: n_3133 <=  gnd;
delay_2601: n_3134  <= TRANSPORT clk  ;
filter_2602: FILTER_a8237

    PORT MAP (IN1 => n_3134, Y => a_SCH1BWORDOUT_F13_G_aCLK);
dff_2603: DFF_a8237

    PORT MAP ( D => a_EQ1040, CLK => a_SCH2BWORDOUT_F13_G_aCLK, CLRN => a_SCH2BWORDOUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F13_G);
inv_2604: a_SCH2BWORDOUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2605: a_EQ1040 <=  n_3143  XOR n_3154;
or3_2606: n_3143 <=  n_3144  OR n_3148  OR n_3151;
and3_2607: n_3144 <=  n_3145  AND n_3146  AND n_3147;
inv_2608: n_3145  <= TRANSPORT NOT a_LC3_D22  ;
inv_2609: n_3146  <= TRANSPORT NOT a_N62_aNOT  ;
delay_2610: n_3147  <= TRANSPORT dbin(5)  ;
and2_2611: n_3148 <=  n_3149  AND n_3150;
delay_2612: n_3149  <= TRANSPORT a_N62_aNOT  ;
delay_2613: n_3150  <= TRANSPORT a_SCH2BWORDOUT_F13_G  ;
and2_2614: n_3151 <=  n_3152  AND n_3153;
delay_2615: n_3152  <= TRANSPORT a_LC3_D22  ;
delay_2616: n_3153  <= TRANSPORT a_SCH2BWORDOUT_F13_G  ;
and1_2617: n_3154 <=  gnd;
delay_2618: n_3155  <= TRANSPORT clk  ;
filter_2619: FILTER_a8237

    PORT MAP (IN1 => n_3155, Y => a_SCH2BWORDOUT_F13_G_aCLK);
dff_2620: DFF_a8237

    PORT MAP ( D => a_EQ1024, CLK => a_SCH2BAROUT_F13_G_aCLK, CLRN => a_SCH2BAROUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F13_G);
inv_2621: a_SCH2BAROUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2622: a_EQ1024 <=  n_3164  XOR n_3171;
or2_2623: n_3164 <=  n_3165  OR n_3168;
and2_2624: n_3165 <=  n_3166  AND n_3167;
inv_2625: n_3166  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_2626: n_3167  <= TRANSPORT dbin(5)  ;
and2_2627: n_3168 <=  n_3169  AND n_3170;
delay_2628: n_3169  <= TRANSPORT a_N2583_aNOT  ;
delay_2629: n_3170  <= TRANSPORT a_SCH2BAROUT_F13_G  ;
and1_2630: n_3171 <=  gnd;
delay_2631: n_3172  <= TRANSPORT clk  ;
filter_2632: FILTER_a8237

    PORT MAP (IN1 => n_3172, Y => a_SCH2BAROUT_F13_G_aCLK);
dff_2633: DFF_a8237

    PORT MAP ( D => a_EQ896, CLK => a_SCH0BAROUT_F13_G_aCLK, CLRN => a_SCH0BAROUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F13_G);
inv_2634: a_SCH0BAROUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2635: a_EQ896 <=  n_3181  XOR n_3188;
or2_2636: n_3181 <=  n_3182  OR n_3185;
and2_2637: n_3182 <=  n_3183  AND n_3184;
inv_2638: n_3183  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_2639: n_3184  <= TRANSPORT dbin(5)  ;
and2_2640: n_3185 <=  n_3186  AND n_3187;
delay_2641: n_3186  <= TRANSPORT a_N2587_aNOT  ;
delay_2642: n_3187  <= TRANSPORT a_SCH0BAROUT_F13_G  ;
and1_2643: n_3188 <=  gnd;
delay_2644: n_3189  <= TRANSPORT clk  ;
filter_2645: FILTER_a8237

    PORT MAP (IN1 => n_3189, Y => a_SCH0BAROUT_F13_G_aCLK);
dff_2646: DFF_a8237

    PORT MAP ( D => a_EQ1088, CLK => a_SCH3BAROUT_F13_G_aCLK, CLRN => a_SCH3BAROUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F13_G);
inv_2647: a_SCH3BAROUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2648: a_EQ1088 <=  n_3198  XOR n_3205;
or2_2649: n_3198 <=  n_3199  OR n_3202;
and2_2650: n_3199 <=  n_3200  AND n_3201;
inv_2651: n_3200  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_2652: n_3201  <= TRANSPORT dbin(5)  ;
and2_2653: n_3202 <=  n_3203  AND n_3204;
delay_2654: n_3203  <= TRANSPORT a_N2581_aNOT  ;
delay_2655: n_3204  <= TRANSPORT a_SCH3BAROUT_F13_G  ;
and1_2656: n_3205 <=  gnd;
delay_2657: n_3206  <= TRANSPORT clk  ;
filter_2658: FILTER_a8237

    PORT MAP (IN1 => n_3206, Y => a_SCH3BAROUT_F13_G_aCLK);
delay_2659: a_LC7_F24  <= TRANSPORT a_EQ807  ;
xor2_2660: a_EQ807 <=  n_3210  XOR n_3220;
or2_2661: n_3210 <=  n_3211  OR n_3215;
and3_2662: n_3211 <=  n_3212  AND n_3213  AND n_3214;
inv_2663: n_3212  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_2664: n_3213  <= TRANSPORT a_N756  ;
delay_2665: n_3214  <= TRANSPORT dbin(6)  ;
and3_2666: n_3215 <=  n_3216  AND n_3217  AND n_3218;
delay_2667: n_3216  <= TRANSPORT a_N2574_aNOT  ;
delay_2668: n_3217  <= TRANSPORT a_N756  ;
delay_2669: n_3218  <= TRANSPORT a_SCH2WRDCNTREG_F6_G  ;
and1_2670: n_3220 <=  gnd;
delay_2671: a_LC7_F13  <= TRANSPORT a_EQ026  ;
xor2_2672: a_EQ026 <=  n_3223  XOR n_3238;
or4_2673: n_3223 <=  n_3224  OR n_3227  OR n_3230  OR n_3233;
and2_2674: n_3224 <=  n_3225  AND n_3226;
delay_2675: n_3225  <= TRANSPORT a_N3552  ;
inv_2676: n_3226  <= TRANSPORT NOT a_N3550  ;
and2_2677: n_3227 <=  n_3228  AND n_3229;
delay_2678: n_3228  <= TRANSPORT a_LC3_C13  ;
inv_2679: n_3229  <= TRANSPORT NOT a_N3550  ;
and2_2680: n_3230 <=  n_3231  AND n_3232;
delay_2681: n_3231  <= TRANSPORT a_N3551  ;
inv_2682: n_3232  <= TRANSPORT NOT a_N3550  ;
and4_2683: n_3233 <=  n_3234  AND n_3235  AND n_3236  AND n_3237;
inv_2684: n_3234  <= TRANSPORT NOT a_LC3_C13  ;
inv_2685: n_3235  <= TRANSPORT NOT a_N3552  ;
inv_2686: n_3236  <= TRANSPORT NOT a_N3551  ;
delay_2687: n_3237  <= TRANSPORT a_N3550  ;
and1_2688: n_3238 <=  gnd;
delay_2689: a_N832_aNOT  <= TRANSPORT a_N832_aNOT_aIN  ;
xor2_2690: a_N832_aNOT_aIN <=  n_3241  XOR n_3246;
or1_2691: n_3241 <=  n_3242;
and3_2692: n_3242 <=  n_3243  AND n_3244  AND n_3245;
inv_2693: n_3243  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_2694: n_3244  <= TRANSPORT NOT a_N2527  ;
inv_2695: n_3245  <= TRANSPORT NOT a_LC7_F13  ;
and1_2696: n_3246 <=  gnd;
dff_2697: DFF_a8237

    PORT MAP ( D => a_EQ1055, CLK => a_SCH2WRDCNTREG_F6_G_aCLK, CLRN => a_SCH2WRDCNTREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F6_G);
inv_2698: a_SCH2WRDCNTREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2699: a_EQ1055 <=  n_3253  XOR n_3261;
or3_2700: n_3253 <=  n_3254  OR n_3256  OR n_3258;
and1_2701: n_3254 <=  n_3255;
delay_2702: n_3255  <= TRANSPORT a_LC7_F24  ;
and1_2703: n_3256 <=  n_3257;
delay_2704: n_3257  <= TRANSPORT a_N832_aNOT  ;
and2_2705: n_3258 <=  n_3259  AND n_3260;
delay_2706: n_3259  <= TRANSPORT a_SCH2BWORDOUT_F6_G  ;
delay_2707: n_3260  <= TRANSPORT a_N2527  ;
and1_2708: n_3261 <=  gnd;
delay_2709: n_3262  <= TRANSPORT clk  ;
filter_2710: FILTER_a8237

    PORT MAP (IN1 => n_3262, Y => a_SCH2WRDCNTREG_F6_G_aCLK);
delay_2711: a_LC5_F27  <= TRANSPORT a_EQ827  ;
xor2_2712: a_EQ827 <=  n_3266  XOR n_3274;
or2_2713: n_3266 <=  n_3267  OR n_3270;
and2_2714: n_3267 <=  n_3268  AND n_3269;
delay_2715: n_3268  <= TRANSPORT a_N1094  ;
inv_2716: n_3269  <= TRANSPORT NOT a_LC7_F13  ;
and2_2717: n_3270 <=  n_3271  AND n_3273;
delay_2718: n_3271  <= TRANSPORT a_SCH3BWORDOUT_F6_G  ;
delay_2719: n_3273  <= TRANSPORT a_N2528  ;
and1_2720: n_3274 <=  gnd;
delay_2721: a_N1066  <= TRANSPORT a_EQ349  ;
xor2_2722: a_EQ349 <=  n_3277  XOR n_3285;
or2_2723: n_3277 <=  n_3278  OR n_3281;
and2_2724: n_3278 <=  n_3279  AND n_3280;
inv_2725: n_3279  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_2726: n_3280  <= TRANSPORT dbin(6)  ;
and2_2727: n_3281 <=  n_3282  AND n_3283;
delay_2728: n_3282  <= TRANSPORT a_N2572_aNOT  ;
delay_2729: n_3283  <= TRANSPORT a_SCH3WRDCNTREG_F6_G  ;
and1_2730: n_3285 <=  gnd;
dff_2731: DFF_a8237

    PORT MAP ( D => a_EQ1119, CLK => a_SCH3WRDCNTREG_F6_G_aCLK, CLRN => a_SCH3WRDCNTREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F6_G);
inv_2732: a_SCH3WRDCNTREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2733: a_EQ1119 <=  n_3292  XOR n_3298;
or2_2734: n_3292 <=  n_3293  OR n_3295;
and1_2735: n_3293 <=  n_3294;
delay_2736: n_3294  <= TRANSPORT a_LC5_F27  ;
and2_2737: n_3295 <=  n_3296  AND n_3297;
delay_2738: n_3296  <= TRANSPORT a_N1095  ;
delay_2739: n_3297  <= TRANSPORT a_N1066  ;
and1_2740: n_3298 <=  gnd;
delay_2741: n_3299  <= TRANSPORT clk  ;
filter_2742: FILTER_a8237

    PORT MAP (IN1 => n_3299, Y => a_SCH3WRDCNTREG_F6_G_aCLK);
delay_2743: a_LC1_F4  <= TRANSPORT a_EQ785  ;
xor2_2744: a_EQ785 <=  n_3303  XOR n_3311;
or2_2745: n_3303 <=  n_3304  OR n_3307;
and2_2746: n_3304 <=  n_3305  AND n_3306;
inv_2747: n_3305  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_2748: n_3306  <= TRANSPORT dbin(6)  ;
and2_2749: n_3307 <=  n_3308  AND n_3309;
delay_2750: n_3308  <= TRANSPORT a_N2576_aNOT  ;
delay_2751: n_3309  <= TRANSPORT a_SCH1WRDCNTREG_F6_G  ;
and1_2752: n_3311 <=  gnd;
delay_2753: a_LC2_F4  <= TRANSPORT a_EQ786  ;
xor2_2754: a_EQ786 <=  n_3314  XOR n_3321;
or2_2755: n_3314 <=  n_3315  OR n_3318;
and2_2756: n_3315 <=  n_3316  AND n_3317;
inv_2757: n_3316  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_2758: n_3317  <= TRANSPORT NOT a_LC7_F13  ;
and2_2759: n_3318 <=  n_3319  AND n_3320;
delay_2760: n_3319  <= TRANSPORT a_N2559_aNOT  ;
delay_2761: n_3320  <= TRANSPORT a_LC1_F4  ;
and1_2762: n_3321 <=  gnd;
dff_2763: DFF_a8237

    PORT MAP ( D => a_EQ991, CLK => a_SCH1WRDCNTREG_F6_G_aCLK, CLRN => a_SCH1WRDCNTREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F6_G);
inv_2764: a_SCH1WRDCNTREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2765: a_EQ991 <=  n_3328  XOR n_3335;
or2_2766: n_3328 <=  n_3329  OR n_3332;
and2_2767: n_3329 <=  n_3330  AND n_3331;
inv_2768: n_3330  <= TRANSPORT NOT a_N2526  ;
delay_2769: n_3331  <= TRANSPORT a_LC2_F4  ;
and2_2770: n_3332 <=  n_3333  AND n_3334;
delay_2771: n_3333  <= TRANSPORT a_SCH1BWORDOUT_F6_G  ;
delay_2772: n_3334  <= TRANSPORT a_N2526  ;
and1_2773: n_3335 <=  gnd;
delay_2774: n_3336  <= TRANSPORT clk  ;
filter_2775: FILTER_a8237

    PORT MAP (IN1 => n_3336, Y => a_SCH1WRDCNTREG_F6_G_aCLK);
delay_2776: a_LC2_F8  <= TRANSPORT a_EQ762  ;
xor2_2777: a_EQ762 <=  n_3340  XOR n_3348;
or2_2778: n_3340 <=  n_3341  OR n_3344;
and2_2779: n_3341 <=  n_3342  AND n_3343;
inv_2780: n_3342  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_2781: n_3343  <= TRANSPORT dbin(6)  ;
and2_2782: n_3344 <=  n_3345  AND n_3346;
delay_2783: n_3345  <= TRANSPORT a_N2578_aNOT  ;
delay_2784: n_3346  <= TRANSPORT a_SCH0WRDCNTREG_F6_G  ;
and1_2785: n_3348 <=  gnd;
delay_2786: a_LC4_F8  <= TRANSPORT a_EQ763  ;
xor2_2787: a_EQ763 <=  n_3351  XOR n_3358;
or2_2788: n_3351 <=  n_3352  OR n_3355;
and2_2789: n_3352 <=  n_3353  AND n_3354;
inv_2790: n_3353  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_2791: n_3354  <= TRANSPORT NOT a_LC7_F13  ;
and2_2792: n_3355 <=  n_3356  AND n_3357;
delay_2793: n_3356  <= TRANSPORT a_N2558_aNOT  ;
delay_2794: n_3357  <= TRANSPORT a_LC2_F8  ;
and1_2795: n_3358 <=  gnd;
dff_2796: DFF_a8237

    PORT MAP ( D => a_EQ927, CLK => a_SCH0WRDCNTREG_F6_G_aCLK, CLRN => a_SCH0WRDCNTREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F6_G);
inv_2797: a_SCH0WRDCNTREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2798: a_EQ927 <=  n_3365  XOR n_3372;
or2_2799: n_3365 <=  n_3366  OR n_3369;
and2_2800: n_3366 <=  n_3367  AND n_3368;
inv_2801: n_3367  <= TRANSPORT NOT a_N2525  ;
delay_2802: n_3368  <= TRANSPORT a_LC4_F8  ;
and2_2803: n_3369 <=  n_3370  AND n_3371;
delay_2804: n_3370  <= TRANSPORT a_SCH0BWORDOUT_F6_G  ;
delay_2805: n_3371  <= TRANSPORT a_N2525  ;
and1_2806: n_3372 <=  gnd;
delay_2807: n_3373  <= TRANSPORT clk  ;
filter_2808: FILTER_a8237

    PORT MAP (IN1 => n_3373, Y => a_SCH0WRDCNTREG_F6_G_aCLK);
dff_2809: DFF_a8237

    PORT MAP ( D => a_EQ897, CLK => a_SCH0BAROUT_F14_G_aCLK, CLRN => a_SCH0BAROUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F14_G);
inv_2810: a_SCH0BAROUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2811: a_EQ897 <=  n_3382  XOR n_3389;
or2_2812: n_3382 <=  n_3383  OR n_3386;
and2_2813: n_3383 <=  n_3384  AND n_3385;
inv_2814: n_3384  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_2815: n_3385  <= TRANSPORT dbin(6)  ;
and2_2816: n_3386 <=  n_3387  AND n_3388;
delay_2817: n_3387  <= TRANSPORT a_N2587_aNOT  ;
delay_2818: n_3388  <= TRANSPORT a_SCH0BAROUT_F14_G  ;
and1_2819: n_3389 <=  gnd;
delay_2820: n_3390  <= TRANSPORT clk  ;
filter_2821: FILTER_a8237

    PORT MAP (IN1 => n_3390, Y => a_SCH0BAROUT_F14_G_aCLK);
dff_2822: DFF_a8237

    PORT MAP ( D => a_EQ1089, CLK => a_SCH3BAROUT_F14_G_aCLK, CLRN => a_SCH3BAROUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F14_G);
inv_2823: a_SCH3BAROUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2824: a_EQ1089 <=  n_3399  XOR n_3406;
or2_2825: n_3399 <=  n_3400  OR n_3403;
and2_2826: n_3400 <=  n_3401  AND n_3402;
inv_2827: n_3401  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_2828: n_3402  <= TRANSPORT dbin(6)  ;
and2_2829: n_3403 <=  n_3404  AND n_3405;
delay_2830: n_3404  <= TRANSPORT a_N2581_aNOT  ;
delay_2831: n_3405  <= TRANSPORT a_SCH3BAROUT_F14_G  ;
and1_2832: n_3406 <=  gnd;
delay_2833: n_3407  <= TRANSPORT clk  ;
filter_2834: FILTER_a8237

    PORT MAP (IN1 => n_3407, Y => a_SCH3BAROUT_F14_G_aCLK);
dff_2835: DFF_a8237

    PORT MAP ( D => a_EQ1098, CLK => a_SCH3BWORDOUT_F7_G_aCLK, CLRN => a_SCH3BWORDOUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F7_G);
inv_2836: a_SCH3BWORDOUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2837: a_EQ1098 <=  n_3416  XOR n_3423;
or2_2838: n_3416 <=  n_3417  OR n_3420;
and2_2839: n_3417 <=  n_3418  AND n_3419;
inv_2840: n_3418  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_2841: n_3419  <= TRANSPORT dbin(7)  ;
and2_2842: n_3420 <=  n_3421  AND n_3422;
delay_2843: n_3421  <= TRANSPORT a_N2572_aNOT  ;
delay_2844: n_3422  <= TRANSPORT a_SCH3BWORDOUT_F7_G  ;
and1_2845: n_3423 <=  gnd;
delay_2846: n_3424  <= TRANSPORT clk  ;
filter_2847: FILTER_a8237

    PORT MAP (IN1 => n_3424, Y => a_SCH3BWORDOUT_F7_G_aCLK);
dff_2848: DFF_a8237

    PORT MAP ( D => a_EQ1034, CLK => a_SCH2BWORDOUT_F7_G_aCLK, CLRN => a_SCH2BWORDOUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F7_G);
inv_2849: a_SCH2BWORDOUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2850: a_EQ1034 <=  n_3433  XOR n_3440;
or2_2851: n_3433 <=  n_3434  OR n_3437;
and2_2852: n_3434 <=  n_3435  AND n_3436;
inv_2853: n_3435  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_2854: n_3436  <= TRANSPORT dbin(7)  ;
and2_2855: n_3437 <=  n_3438  AND n_3439;
delay_2856: n_3438  <= TRANSPORT a_N2574_aNOT  ;
delay_2857: n_3439  <= TRANSPORT a_SCH2BWORDOUT_F7_G  ;
and1_2858: n_3440 <=  gnd;
delay_2859: n_3441  <= TRANSPORT clk  ;
filter_2860: FILTER_a8237

    PORT MAP (IN1 => n_3441, Y => a_SCH2BWORDOUT_F7_G_aCLK);
dff_2861: DFF_a8237

    PORT MAP ( D => a_EQ906, CLK => a_SCH0BWORDOUT_F7_G_aCLK, CLRN => a_SCH0BWORDOUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F7_G);
inv_2862: a_SCH0BWORDOUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2863: a_EQ906 <=  n_3450  XOR n_3457;
or2_2864: n_3450 <=  n_3451  OR n_3454;
and2_2865: n_3451 <=  n_3452  AND n_3453;
inv_2866: n_3452  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_2867: n_3453  <= TRANSPORT dbin(7)  ;
and2_2868: n_3454 <=  n_3455  AND n_3456;
delay_2869: n_3455  <= TRANSPORT a_N2578_aNOT  ;
delay_2870: n_3456  <= TRANSPORT a_SCH0BWORDOUT_F7_G  ;
and1_2871: n_3457 <=  gnd;
delay_2872: n_3458  <= TRANSPORT clk  ;
filter_2873: FILTER_a8237

    PORT MAP (IN1 => n_3458, Y => a_SCH0BWORDOUT_F7_G_aCLK);
dff_2874: DFF_a8237

    PORT MAP ( D => a_EQ1026, CLK => a_SCH2BAROUT_F15_G_aCLK, CLRN => a_SCH2BAROUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F15_G);
inv_2875: a_SCH2BAROUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2876: a_EQ1026 <=  n_3467  XOR n_3474;
or2_2877: n_3467 <=  n_3468  OR n_3471;
and2_2878: n_3468 <=  n_3469  AND n_3470;
inv_2879: n_3469  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_2880: n_3470  <= TRANSPORT dbin(7)  ;
and2_2881: n_3471 <=  n_3472  AND n_3473;
delay_2882: n_3472  <= TRANSPORT a_N2583_aNOT  ;
delay_2883: n_3473  <= TRANSPORT a_SCH2BAROUT_F15_G  ;
and1_2884: n_3474 <=  gnd;
delay_2885: n_3475  <= TRANSPORT clk  ;
filter_2886: FILTER_a8237

    PORT MAP (IN1 => n_3475, Y => a_SCH2BAROUT_F15_G_aCLK);
dff_2887: DFF_a8237

    PORT MAP ( D => a_EQ898, CLK => a_SCH0BAROUT_F15_G_aCLK, CLRN => a_SCH0BAROUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F15_G);
inv_2888: a_SCH0BAROUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2889: a_EQ898 <=  n_3484  XOR n_3491;
or2_2890: n_3484 <=  n_3485  OR n_3488;
and2_2891: n_3485 <=  n_3486  AND n_3487;
delay_2892: n_3486  <= TRANSPORT a_N2587_aNOT  ;
delay_2893: n_3487  <= TRANSPORT a_SCH0BAROUT_F15_G  ;
and2_2894: n_3488 <=  n_3489  AND n_3490;
inv_2895: n_3489  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_2896: n_3490  <= TRANSPORT dbin(7)  ;
and1_2897: n_3491 <=  gnd;
delay_2898: n_3492  <= TRANSPORT clk  ;
filter_2899: FILTER_a8237

    PORT MAP (IN1 => n_3492, Y => a_SCH0BAROUT_F15_G_aCLK);
dff_2900: DFF_a8237

    PORT MAP ( D => a_EQ1090, CLK => a_SCH3BAROUT_F15_G_aCLK, CLRN => a_SCH3BAROUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F15_G);
inv_2901: a_SCH3BAROUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2902: a_EQ1090 <=  n_3501  XOR n_3508;
or2_2903: n_3501 <=  n_3502  OR n_3505;
and2_2904: n_3502 <=  n_3503  AND n_3504;
inv_2905: n_3503  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_2906: n_3504  <= TRANSPORT dbin(7)  ;
and2_2907: n_3505 <=  n_3506  AND n_3507;
delay_2908: n_3506  <= TRANSPORT a_N2581_aNOT  ;
delay_2909: n_3507  <= TRANSPORT a_SCH3BAROUT_F15_G  ;
and1_2910: n_3508 <=  gnd;
delay_2911: n_3509  <= TRANSPORT clk  ;
filter_2912: FILTER_a8237

    PORT MAP (IN1 => n_3509, Y => a_SCH3BAROUT_F15_G_aCLK);
dff_2913: DFF_a8237

    PORT MAP ( D => a_EQ962, CLK => a_SCH1BAROUT_F15_G_aCLK, CLRN => a_SCH1BAROUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F15_G);
inv_2914: a_SCH1BAROUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2915: a_EQ962 <=  n_3518  XOR n_3525;
or2_2916: n_3518 <=  n_3519  OR n_3522;
and2_2917: n_3519 <=  n_3520  AND n_3521;
inv_2918: n_3520  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_2919: n_3521  <= TRANSPORT dbin(7)  ;
and2_2920: n_3522 <=  n_3523  AND n_3524;
delay_2921: n_3523  <= TRANSPORT a_N2585_aNOT  ;
delay_2922: n_3524  <= TRANSPORT a_SCH1BAROUT_F15_G  ;
and1_2923: n_3525 <=  gnd;
delay_2924: n_3526  <= TRANSPORT clk  ;
filter_2925: FILTER_a8237

    PORT MAP (IN1 => n_3526, Y => a_SCH1BAROUT_F15_G_aCLK);
delay_2926: a_LC5_A20  <= TRANSPORT a_EQ029  ;
xor2_2927: a_EQ029 <=  n_3530  XOR n_3541;
or3_2928: n_3530 <=  n_3531  OR n_3534  OR n_3537;
and2_2929: n_3531 <=  n_3532  AND n_3533;
delay_2930: n_3532  <= TRANSPORT a_N3546  ;
inv_2931: n_3533  <= TRANSPORT NOT a_N3545  ;
and2_2932: n_3534 <=  n_3535  AND n_3536;
inv_2933: n_3535  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
inv_2934: n_3536  <= TRANSPORT NOT a_N3545  ;
and3_2935: n_3537 <=  n_3538  AND n_3539  AND n_3540;
delay_2936: n_3538  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_2937: n_3539  <= TRANSPORT NOT a_N3546  ;
delay_2938: n_3540  <= TRANSPORT a_N3545  ;
and1_2939: n_3541 <=  gnd;
delay_2940: a_LC4_A22  <= TRANSPORT a_EQ820  ;
xor2_2941: a_EQ820 <=  n_3544  XOR n_3552;
or2_2942: n_3544 <=  n_3545  OR n_3548;
and2_2943: n_3545 <=  n_3546  AND n_3547;
inv_2944: n_3546  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_2945: n_3547  <= TRANSPORT dbin(3)  ;
and2_2946: n_3548 <=  n_3549  AND n_3550;
delay_2947: n_3549  <= TRANSPORT a_N2573_aNOT  ;
delay_2948: n_3550  <= TRANSPORT a_SH3WRDCNTREG_F11_G  ;
and1_2949: n_3552 <=  gnd;
delay_2950: a_LC3_A22  <= TRANSPORT a_EQ821  ;
xor2_2951: a_EQ821 <=  n_3555  XOR n_3562;
or2_2952: n_3555 <=  n_3556  OR n_3559;
and2_2953: n_3556 <=  n_3557  AND n_3558;
inv_2954: n_3557  <= TRANSPORT NOT a_N965  ;
inv_2955: n_3558  <= TRANSPORT NOT a_LC5_A20  ;
and2_2956: n_3559 <=  n_3560  AND n_3561;
delay_2957: n_3560  <= TRANSPORT a_N965  ;
delay_2958: n_3561  <= TRANSPORT a_LC4_A22  ;
and1_2959: n_3562 <=  gnd;
dff_2960: DFF_a8237

    PORT MAP ( D => a_EQ1152, CLK => a_SH3WRDCNTREG_F11_G_aCLK, CLRN => a_SH3WRDCNTREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SH3WRDCNTREG_F11_G);
inv_2961: a_SH3WRDCNTREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2962: a_EQ1152 <=  n_3569  XOR n_3576;
or2_2963: n_3569 <=  n_3570  OR n_3573;
and2_2964: n_3570 <=  n_3571  AND n_3572;
inv_2965: n_3571  <= TRANSPORT NOT a_N2528  ;
delay_2966: n_3572  <= TRANSPORT a_LC3_A22  ;
and2_2967: n_3573 <=  n_3574  AND n_3575;
delay_2968: n_3574  <= TRANSPORT a_SCH3BWORDOUT_F11_G  ;
delay_2969: n_3575  <= TRANSPORT a_N2528  ;
and1_2970: n_3576 <=  gnd;
delay_2971: n_3577  <= TRANSPORT clk  ;
filter_2972: FILTER_a8237

    PORT MAP (IN1 => n_3577, Y => a_SH3WRDCNTREG_F11_G_aCLK);
delay_2973: a_LC5_A11  <= TRANSPORT a_EQ778  ;
xor2_2974: a_EQ778 <=  n_3581  XOR n_3589;
or2_2975: n_3581 <=  n_3582  OR n_3585;
and2_2976: n_3582 <=  n_3583  AND n_3584;
inv_2977: n_3583  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_2978: n_3584  <= TRANSPORT dbin(3)  ;
and2_2979: n_3585 <=  n_3586  AND n_3587;
delay_2980: n_3586  <= TRANSPORT a_N2577_aNOT  ;
delay_2981: n_3587  <= TRANSPORT a_SH1WRDCNTREG_F11_G  ;
and1_2982: n_3589 <=  gnd;
delay_2983: a_LC3_A11  <= TRANSPORT a_EQ779  ;
xor2_2984: a_EQ779 <=  n_3592  XOR n_3599;
or2_2985: n_3592 <=  n_3593  OR n_3596;
and2_2986: n_3593 <=  n_3594  AND n_3595;
inv_2987: n_3594  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_2988: n_3595  <= TRANSPORT NOT a_LC5_A20  ;
and2_2989: n_3596 <=  n_3597  AND n_3598;
delay_2990: n_3597  <= TRANSPORT a_N2559_aNOT  ;
delay_2991: n_3598  <= TRANSPORT a_LC5_A11  ;
and1_2992: n_3599 <=  gnd;
dff_2993: DFF_a8237

    PORT MAP ( D => a_EQ1140, CLK => a_SH1WRDCNTREG_F11_G_aCLK, CLRN => a_SH1WRDCNTREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SH1WRDCNTREG_F11_G);
inv_2994: a_SH1WRDCNTREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_2995: a_EQ1140 <=  n_3606  XOR n_3613;
or2_2996: n_3606 <=  n_3607  OR n_3610;
and2_2997: n_3607 <=  n_3608  AND n_3609;
inv_2998: n_3608  <= TRANSPORT NOT a_N2526  ;
delay_2999: n_3609  <= TRANSPORT a_LC3_A11  ;
and2_3000: n_3610 <=  n_3611  AND n_3612;
delay_3001: n_3611  <= TRANSPORT a_SCH1BWORDOUT_F11_G  ;
delay_3002: n_3612  <= TRANSPORT a_N2526  ;
and1_3003: n_3613 <=  gnd;
delay_3004: n_3614  <= TRANSPORT clk  ;
filter_3005: FILTER_a8237

    PORT MAP (IN1 => n_3614, Y => a_SH1WRDCNTREG_F11_G_aCLK);
delay_3006: a_LC4_F26  <= TRANSPORT a_EQ799  ;
xor2_3007: a_EQ799 <=  n_3618  XOR n_3630;
or3_3008: n_3618 <=  n_3619  OR n_3623  OR n_3627;
and3_3009: n_3619 <=  n_3620  AND n_3621  AND n_3622;
inv_3010: n_3620  <= TRANSPORT NOT a_LC3_D22  ;
inv_3011: n_3621  <= TRANSPORT NOT a_N62_aNOT  ;
delay_3012: n_3622  <= TRANSPORT dbin(3)  ;
and2_3013: n_3623 <=  n_3624  AND n_3625;
delay_3014: n_3624  <= TRANSPORT a_N62_aNOT  ;
delay_3015: n_3625  <= TRANSPORT a_SH2WRDCNTREG_F11_G  ;
and2_3016: n_3627 <=  n_3628  AND n_3629;
delay_3017: n_3628  <= TRANSPORT a_LC3_D22  ;
delay_3018: n_3629  <= TRANSPORT a_SH2WRDCNTREG_F11_G  ;
and1_3019: n_3630 <=  gnd;
delay_3020: a_LC5_F26  <= TRANSPORT a_EQ800  ;
xor2_3021: a_EQ800 <=  n_3633  XOR n_3640;
or2_3022: n_3633 <=  n_3634  OR n_3637;
and2_3023: n_3634 <=  n_3635  AND n_3636;
inv_3024: n_3635  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_3025: n_3636  <= TRANSPORT NOT a_LC5_A20  ;
and2_3026: n_3637 <=  n_3638  AND n_3639;
delay_3027: n_3638  <= TRANSPORT a_N2560_aNOT  ;
delay_3028: n_3639  <= TRANSPORT a_LC4_F26  ;
and1_3029: n_3640 <=  gnd;
dff_3030: DFF_a8237

    PORT MAP ( D => a_EQ1146, CLK => a_SH2WRDCNTREG_F11_G_aCLK, CLRN => a_SH2WRDCNTREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SH2WRDCNTREG_F11_G);
inv_3031: a_SH2WRDCNTREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3032: a_EQ1146 <=  n_3647  XOR n_3654;
or2_3033: n_3647 <=  n_3648  OR n_3651;
and2_3034: n_3648 <=  n_3649  AND n_3650;
inv_3035: n_3649  <= TRANSPORT NOT a_N2527  ;
delay_3036: n_3650  <= TRANSPORT a_LC5_F26  ;
and2_3037: n_3651 <=  n_3652  AND n_3653;
delay_3038: n_3652  <= TRANSPORT a_SCH2BWORDOUT_F11_G  ;
delay_3039: n_3653  <= TRANSPORT a_N2527  ;
and1_3040: n_3654 <=  gnd;
delay_3041: n_3655  <= TRANSPORT clk  ;
filter_3042: FILTER_a8237

    PORT MAP (IN1 => n_3655, Y => a_SH2WRDCNTREG_F11_G_aCLK);
delay_3043: a_LC5_A22  <= TRANSPORT a_EQ756  ;
xor2_3044: a_EQ756 <=  n_3659  XOR n_3671;
or3_3045: n_3659 <=  n_3660  OR n_3664  OR n_3668;
and3_3046: n_3660 <=  n_3661  AND n_3662  AND n_3663;
inv_3047: n_3661  <= TRANSPORT NOT a_LC3_D22  ;
inv_3048: n_3662  <= TRANSPORT NOT a_N2353  ;
delay_3049: n_3663  <= TRANSPORT dbin(3)  ;
and2_3050: n_3664 <=  n_3665  AND n_3666;
delay_3051: n_3665  <= TRANSPORT a_N2353  ;
delay_3052: n_3666  <= TRANSPORT a_SH0WRDCNTREG_F11_G  ;
and2_3053: n_3668 <=  n_3669  AND n_3670;
delay_3054: n_3669  <= TRANSPORT a_LC3_D22  ;
delay_3055: n_3670  <= TRANSPORT a_SH0WRDCNTREG_F11_G  ;
and1_3056: n_3671 <=  gnd;
delay_3057: a_LC6_A22  <= TRANSPORT a_EQ757  ;
xor2_3058: a_EQ757 <=  n_3674  XOR n_3681;
or2_3059: n_3674 <=  n_3675  OR n_3678;
and2_3060: n_3675 <=  n_3676  AND n_3677;
inv_3061: n_3676  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_3062: n_3677  <= TRANSPORT NOT a_LC5_A20  ;
and2_3063: n_3678 <=  n_3679  AND n_3680;
delay_3064: n_3679  <= TRANSPORT a_N2558_aNOT  ;
delay_3065: n_3680  <= TRANSPORT a_LC5_A22  ;
and1_3066: n_3681 <=  gnd;
dff_3067: DFF_a8237

    PORT MAP ( D => a_EQ1134, CLK => a_SH0WRDCNTREG_F11_G_aCLK, CLRN => a_SH0WRDCNTREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SH0WRDCNTREG_F11_G);
inv_3068: a_SH0WRDCNTREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3069: a_EQ1134 <=  n_3688  XOR n_3695;
or2_3070: n_3688 <=  n_3689  OR n_3692;
and2_3071: n_3689 <=  n_3690  AND n_3691;
inv_3072: n_3690  <= TRANSPORT NOT a_N2525  ;
delay_3073: n_3691  <= TRANSPORT a_LC6_A22  ;
and2_3074: n_3692 <=  n_3693  AND n_3694;
delay_3075: n_3693  <= TRANSPORT a_SCH0BWORDOUT_F11_G  ;
delay_3076: n_3694  <= TRANSPORT a_N2525  ;
and1_3077: n_3695 <=  gnd;
delay_3078: n_3696  <= TRANSPORT clk  ;
filter_3079: FILTER_a8237

    PORT MAP (IN1 => n_3696, Y => a_SH0WRDCNTREG_F11_G_aCLK);
delay_3080: a_LC6_A20  <= TRANSPORT a_EQ030  ;
xor2_3081: a_EQ030 <=  n_3700  XOR n_3715;
or4_3082: n_3700 <=  n_3701  OR n_3704  OR n_3707  OR n_3710;
and2_3083: n_3701 <=  n_3702  AND n_3703;
delay_3084: n_3702  <= TRANSPORT a_N3545  ;
inv_3085: n_3703  <= TRANSPORT NOT a_N3544  ;
and2_3086: n_3704 <=  n_3705  AND n_3706;
delay_3087: n_3705  <= TRANSPORT a_N3546  ;
inv_3088: n_3706  <= TRANSPORT NOT a_N3544  ;
and2_3089: n_3707 <=  n_3708  AND n_3709;
inv_3090: n_3708  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
inv_3091: n_3709  <= TRANSPORT NOT a_N3544  ;
and4_3092: n_3710 <=  n_3711  AND n_3712  AND n_3713  AND n_3714;
delay_3093: n_3711  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_3094: n_3712  <= TRANSPORT NOT a_N3546  ;
inv_3095: n_3713  <= TRANSPORT NOT a_N3545  ;
delay_3096: n_3714  <= TRANSPORT a_N3544  ;
and1_3097: n_3715 <=  gnd;
delay_3098: a_LC3_A21  <= TRANSPORT a_EQ818  ;
xor2_3099: a_EQ818 <=  n_3718  XOR n_3726;
or2_3100: n_3718 <=  n_3719  OR n_3722;
and2_3101: n_3719 <=  n_3720  AND n_3721;
inv_3102: n_3720  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_3103: n_3721  <= TRANSPORT dbin(4)  ;
and2_3104: n_3722 <=  n_3723  AND n_3724;
delay_3105: n_3723  <= TRANSPORT a_N2573_aNOT  ;
delay_3106: n_3724  <= TRANSPORT a_SH3WRDCNTREG_F12_G  ;
and1_3107: n_3726 <=  gnd;
delay_3108: a_LC4_A21  <= TRANSPORT a_EQ819  ;
xor2_3109: a_EQ819 <=  n_3729  XOR n_3736;
or2_3110: n_3729 <=  n_3730  OR n_3733;
and2_3111: n_3730 <=  n_3731  AND n_3732;
inv_3112: n_3731  <= TRANSPORT NOT a_N965  ;
inv_3113: n_3732  <= TRANSPORT NOT a_LC6_A20  ;
and2_3114: n_3733 <=  n_3734  AND n_3735;
delay_3115: n_3734  <= TRANSPORT a_N965  ;
delay_3116: n_3735  <= TRANSPORT a_LC3_A21  ;
and1_3117: n_3736 <=  gnd;
dff_3118: DFF_a8237

    PORT MAP ( D => a_EQ1153, CLK => a_SH3WRDCNTREG_F12_G_aCLK, CLRN => a_SH3WRDCNTREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SH3WRDCNTREG_F12_G);
inv_3119: a_SH3WRDCNTREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3120: a_EQ1153 <=  n_3743  XOR n_3750;
or2_3121: n_3743 <=  n_3744  OR n_3747;
and2_3122: n_3744 <=  n_3745  AND n_3746;
inv_3123: n_3745  <= TRANSPORT NOT a_N2528  ;
delay_3124: n_3746  <= TRANSPORT a_LC4_A21  ;
and2_3125: n_3747 <=  n_3748  AND n_3749;
delay_3126: n_3748  <= TRANSPORT a_SCH3BWORDOUT_F12_G  ;
delay_3127: n_3749  <= TRANSPORT a_N2528  ;
and1_3128: n_3750 <=  gnd;
delay_3129: n_3751  <= TRANSPORT clk  ;
filter_3130: FILTER_a8237

    PORT MAP (IN1 => n_3751, Y => a_SH3WRDCNTREG_F12_G_aCLK);
delay_3131: a_LC1_A8  <= TRANSPORT a_EQ754  ;
xor2_3132: a_EQ754 <=  n_3755  XOR n_3767;
or3_3133: n_3755 <=  n_3756  OR n_3760  OR n_3764;
and3_3134: n_3756 <=  n_3757  AND n_3758  AND n_3759;
inv_3135: n_3757  <= TRANSPORT NOT a_LC3_D22  ;
inv_3136: n_3758  <= TRANSPORT NOT a_N2353  ;
delay_3137: n_3759  <= TRANSPORT dbin(4)  ;
and2_3138: n_3760 <=  n_3761  AND n_3762;
delay_3139: n_3761  <= TRANSPORT a_N2353  ;
delay_3140: n_3762  <= TRANSPORT a_SH0WRDCNTREG_F12_G  ;
and2_3141: n_3764 <=  n_3765  AND n_3766;
delay_3142: n_3765  <= TRANSPORT a_LC3_D22  ;
delay_3143: n_3766  <= TRANSPORT a_SH0WRDCNTREG_F12_G  ;
and1_3144: n_3767 <=  gnd;
delay_3145: a_LC2_A8  <= TRANSPORT a_EQ755  ;
xor2_3146: a_EQ755 <=  n_3770  XOR n_3777;
or2_3147: n_3770 <=  n_3771  OR n_3774;
and2_3148: n_3771 <=  n_3772  AND n_3773;
inv_3149: n_3772  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_3150: n_3773  <= TRANSPORT NOT a_LC6_A20  ;
and2_3151: n_3774 <=  n_3775  AND n_3776;
delay_3152: n_3775  <= TRANSPORT a_N2558_aNOT  ;
delay_3153: n_3776  <= TRANSPORT a_LC1_A8  ;
and1_3154: n_3777 <=  gnd;
dff_3155: DFF_a8237

    PORT MAP ( D => a_EQ1135, CLK => a_SH0WRDCNTREG_F12_G_aCLK, CLRN => a_SH0WRDCNTREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SH0WRDCNTREG_F12_G);
inv_3156: a_SH0WRDCNTREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3157: a_EQ1135 <=  n_3784  XOR n_3791;
or2_3158: n_3784 <=  n_3785  OR n_3788;
and2_3159: n_3785 <=  n_3786  AND n_3787;
inv_3160: n_3786  <= TRANSPORT NOT a_N2525  ;
delay_3161: n_3787  <= TRANSPORT a_LC2_A8  ;
and2_3162: n_3788 <=  n_3789  AND n_3790;
delay_3163: n_3789  <= TRANSPORT a_SCH0BWORDOUT_F12_G  ;
delay_3164: n_3790  <= TRANSPORT a_N2525  ;
and1_3165: n_3791 <=  gnd;
delay_3166: n_3792  <= TRANSPORT clk  ;
filter_3167: FILTER_a8237

    PORT MAP (IN1 => n_3792, Y => a_SH0WRDCNTREG_F12_G_aCLK);
delay_3168: a_LC3_A14  <= TRANSPORT a_EQ797  ;
xor2_3169: a_EQ797 <=  n_3796  XOR n_3808;
or3_3170: n_3796 <=  n_3797  OR n_3801  OR n_3805;
and3_3171: n_3797 <=  n_3798  AND n_3799  AND n_3800;
inv_3172: n_3798  <= TRANSPORT NOT a_LC3_D22  ;
inv_3173: n_3799  <= TRANSPORT NOT a_N62_aNOT  ;
delay_3174: n_3800  <= TRANSPORT dbin(4)  ;
and2_3175: n_3801 <=  n_3802  AND n_3803;
delay_3176: n_3802  <= TRANSPORT a_N62_aNOT  ;
delay_3177: n_3803  <= TRANSPORT a_SH2WRDCNTREG_F12_G  ;
and2_3178: n_3805 <=  n_3806  AND n_3807;
delay_3179: n_3806  <= TRANSPORT a_LC3_D22  ;
delay_3180: n_3807  <= TRANSPORT a_SH2WRDCNTREG_F12_G  ;
and1_3181: n_3808 <=  gnd;
delay_3182: a_LC2_A14  <= TRANSPORT a_EQ798  ;
xor2_3183: a_EQ798 <=  n_3811  XOR n_3818;
or2_3184: n_3811 <=  n_3812  OR n_3815;
and2_3185: n_3812 <=  n_3813  AND n_3814;
inv_3186: n_3813  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_3187: n_3814  <= TRANSPORT NOT a_LC6_A20  ;
and2_3188: n_3815 <=  n_3816  AND n_3817;
delay_3189: n_3816  <= TRANSPORT a_N2560_aNOT  ;
delay_3190: n_3817  <= TRANSPORT a_LC3_A14  ;
and1_3191: n_3818 <=  gnd;
dff_3192: DFF_a8237

    PORT MAP ( D => a_EQ1147, CLK => a_SH2WRDCNTREG_F12_G_aCLK, CLRN => a_SH2WRDCNTREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SH2WRDCNTREG_F12_G);
inv_3193: a_SH2WRDCNTREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3194: a_EQ1147 <=  n_3825  XOR n_3832;
or2_3195: n_3825 <=  n_3826  OR n_3829;
and2_3196: n_3826 <=  n_3827  AND n_3828;
inv_3197: n_3827  <= TRANSPORT NOT a_N2527  ;
delay_3198: n_3828  <= TRANSPORT a_LC2_A14  ;
and2_3199: n_3829 <=  n_3830  AND n_3831;
delay_3200: n_3830  <= TRANSPORT a_SCH2BWORDOUT_F12_G  ;
delay_3201: n_3831  <= TRANSPORT a_N2527  ;
and1_3202: n_3832 <=  gnd;
delay_3203: n_3833  <= TRANSPORT clk  ;
filter_3204: FILTER_a8237

    PORT MAP (IN1 => n_3833, Y => a_SH2WRDCNTREG_F12_G_aCLK);
delay_3205: a_LC1_A11  <= TRANSPORT a_EQ776  ;
xor2_3206: a_EQ776 <=  n_3837  XOR n_3845;
or2_3207: n_3837 <=  n_3838  OR n_3841;
and2_3208: n_3838 <=  n_3839  AND n_3840;
inv_3209: n_3839  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_3210: n_3840  <= TRANSPORT dbin(4)  ;
and2_3211: n_3841 <=  n_3842  AND n_3843;
delay_3212: n_3842  <= TRANSPORT a_N2577_aNOT  ;
delay_3213: n_3843  <= TRANSPORT a_SH1WRDCNTREG_F12_G  ;
and1_3214: n_3845 <=  gnd;
delay_3215: a_LC2_A11  <= TRANSPORT a_EQ777  ;
xor2_3216: a_EQ777 <=  n_3848  XOR n_3855;
or2_3217: n_3848 <=  n_3849  OR n_3852;
and2_3218: n_3849 <=  n_3850  AND n_3851;
inv_3219: n_3850  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_3220: n_3851  <= TRANSPORT NOT a_LC6_A20  ;
and2_3221: n_3852 <=  n_3853  AND n_3854;
delay_3222: n_3853  <= TRANSPORT a_N2559_aNOT  ;
delay_3223: n_3854  <= TRANSPORT a_LC1_A11  ;
and1_3224: n_3855 <=  gnd;
dff_3225: DFF_a8237

    PORT MAP ( D => a_EQ1141, CLK => a_SH1WRDCNTREG_F12_G_aCLK, CLRN => a_SH1WRDCNTREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SH1WRDCNTREG_F12_G);
inv_3226: a_SH1WRDCNTREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3227: a_EQ1141 <=  n_3862  XOR n_3869;
or2_3228: n_3862 <=  n_3863  OR n_3866;
and2_3229: n_3863 <=  n_3864  AND n_3865;
inv_3230: n_3864  <= TRANSPORT NOT a_N2526  ;
delay_3231: n_3865  <= TRANSPORT a_LC2_A11  ;
and2_3232: n_3866 <=  n_3867  AND n_3868;
delay_3233: n_3867  <= TRANSPORT a_SCH1BWORDOUT_F12_G  ;
delay_3234: n_3868  <= TRANSPORT a_N2526  ;
and1_3235: n_3869 <=  gnd;
delay_3236: n_3870  <= TRANSPORT clk  ;
filter_3237: FILTER_a8237

    PORT MAP (IN1 => n_3870, Y => a_SH1WRDCNTREG_F12_G_aCLK);
dff_3238: DFF_a8237

    PORT MAP ( D => a_EQ914, CLK => a_SCH0BWORDOUT_F15_G_aCLK, CLRN => a_SCH0BWORDOUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F15_G);
inv_3239: a_SCH0BWORDOUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3240: a_EQ914 <=  n_3879  XOR n_3890;
or3_3241: n_3879 <=  n_3880  OR n_3884  OR n_3887;
and3_3242: n_3880 <=  n_3881  AND n_3882  AND n_3883;
inv_3243: n_3881  <= TRANSPORT NOT a_LC3_D22  ;
inv_3244: n_3882  <= TRANSPORT NOT a_N2353  ;
delay_3245: n_3883  <= TRANSPORT dbin(7)  ;
and2_3246: n_3884 <=  n_3885  AND n_3886;
delay_3247: n_3885  <= TRANSPORT a_N2353  ;
delay_3248: n_3886  <= TRANSPORT a_SCH0BWORDOUT_F15_G  ;
and2_3249: n_3887 <=  n_3888  AND n_3889;
delay_3250: n_3888  <= TRANSPORT a_LC3_D22  ;
delay_3251: n_3889  <= TRANSPORT a_SCH0BWORDOUT_F15_G  ;
and1_3252: n_3890 <=  gnd;
delay_3253: n_3891  <= TRANSPORT clk  ;
filter_3254: FILTER_a8237

    PORT MAP (IN1 => n_3891, Y => a_SCH0BWORDOUT_F15_G_aCLK);
dff_3255: DFF_a8237

    PORT MAP ( D => a_EQ978, CLK => a_SCH1BWORDOUT_F15_G_aCLK, CLRN => a_SCH1BWORDOUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F15_G);
inv_3256: a_SCH1BWORDOUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3257: a_EQ978 <=  n_3900  XOR n_3907;
or2_3258: n_3900 <=  n_3901  OR n_3904;
and2_3259: n_3901 <=  n_3902  AND n_3903;
inv_3260: n_3902  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_3261: n_3903  <= TRANSPORT dbin(7)  ;
and2_3262: n_3904 <=  n_3905  AND n_3906;
delay_3263: n_3905  <= TRANSPORT a_N2577_aNOT  ;
delay_3264: n_3906  <= TRANSPORT a_SCH1BWORDOUT_F15_G  ;
and1_3265: n_3907 <=  gnd;
delay_3266: n_3908  <= TRANSPORT clk  ;
filter_3267: FILTER_a8237

    PORT MAP (IN1 => n_3908, Y => a_SCH1BWORDOUT_F15_G_aCLK);
dff_3268: DFF_a8237

    PORT MAP ( D => a_EQ1042, CLK => a_SCH2BWORDOUT_F15_G_aCLK, CLRN => a_SCH2BWORDOUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F15_G);
inv_3269: a_SCH2BWORDOUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3270: a_EQ1042 <=  n_3917  XOR n_3928;
or3_3271: n_3917 <=  n_3918  OR n_3922  OR n_3925;
and3_3272: n_3918 <=  n_3919  AND n_3920  AND n_3921;
inv_3273: n_3919  <= TRANSPORT NOT a_LC3_D22  ;
inv_3274: n_3920  <= TRANSPORT NOT a_N62_aNOT  ;
delay_3275: n_3921  <= TRANSPORT dbin(7)  ;
and2_3276: n_3922 <=  n_3923  AND n_3924;
delay_3277: n_3923  <= TRANSPORT a_N62_aNOT  ;
delay_3278: n_3924  <= TRANSPORT a_SCH2BWORDOUT_F15_G  ;
and2_3279: n_3925 <=  n_3926  AND n_3927;
delay_3280: n_3926  <= TRANSPORT a_LC3_D22  ;
delay_3281: n_3927  <= TRANSPORT a_SCH2BWORDOUT_F15_G  ;
and1_3282: n_3928 <=  gnd;
delay_3283: n_3929  <= TRANSPORT clk  ;
filter_3284: FILTER_a8237

    PORT MAP (IN1 => n_3929, Y => a_SCH2BWORDOUT_F15_G_aCLK);
dff_3285: DFF_a8237

    PORT MAP ( D => a_EQ1106, CLK => a_SCH3BWORDOUT_F15_G_aCLK, CLRN => a_SCH3BWORDOUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F15_G);
inv_3286: a_SCH3BWORDOUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3287: a_EQ1106 <=  n_3938  XOR n_3945;
or2_3288: n_3938 <=  n_3939  OR n_3942;
and2_3289: n_3939 <=  n_3940  AND n_3941;
inv_3290: n_3940  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_3291: n_3941  <= TRANSPORT dbin(7)  ;
and2_3292: n_3942 <=  n_3943  AND n_3944;
delay_3293: n_3943  <= TRANSPORT a_N2573_aNOT  ;
delay_3294: n_3944  <= TRANSPORT a_SCH3BWORDOUT_F15_G  ;
and1_3295: n_3945 <=  gnd;
delay_3296: n_3946  <= TRANSPORT clk  ;
filter_3297: FILTER_a8237

    PORT MAP (IN1 => n_3946, Y => a_SCH3BWORDOUT_F15_G_aCLK);
delay_3298: a_LC6_E16  <= TRANSPORT a_EQ031  ;
xor2_3299: a_EQ031 <=  n_3950  XOR n_3961;
or3_3300: n_3950 <=  n_3951  OR n_3954  OR n_3957;
and2_3301: n_3951 <=  n_3952  AND n_3953;
delay_3302: n_3952  <= TRANSPORT a_N3543  ;
inv_3303: n_3953  <= TRANSPORT NOT a_N3542  ;
and2_3304: n_3954 <=  n_3955  AND n_3956;
inv_3305: n_3955  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
inv_3306: n_3956  <= TRANSPORT NOT a_N3542  ;
and3_3307: n_3957 <=  n_3958  AND n_3959  AND n_3960;
delay_3308: n_3958  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_3309: n_3959  <= TRANSPORT NOT a_N3543  ;
delay_3310: n_3960  <= TRANSPORT a_N3542  ;
and1_3311: n_3961 <=  gnd;
delay_3312: a_LC6_E5  <= TRANSPORT a_EQ352  ;
xor2_3313: a_EQ352 <=  n_3964  XOR n_3972;
or2_3314: n_3964 <=  n_3965  OR n_3968;
and2_3315: n_3965 <=  n_3966  AND n_3967;
inv_3316: n_3966  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_3317: n_3967  <= TRANSPORT dbin(6)  ;
and2_3318: n_3968 <=  n_3969  AND n_3970;
delay_3319: n_3969  <= TRANSPORT a_N2573_aNOT  ;
delay_3320: n_3970  <= TRANSPORT a_SH3WRDCNTREG_F14_G  ;
and1_3321: n_3972 <=  gnd;
delay_3322: a_LC5_E5  <= TRANSPORT a_EQ646  ;
xor2_3323: a_EQ646 <=  n_3975  XOR n_3982;
or2_3324: n_3975 <=  n_3976  OR n_3979;
and2_3325: n_3976 <=  n_3977  AND n_3978;
inv_3326: n_3977  <= TRANSPORT NOT a_N965  ;
inv_3327: n_3978  <= TRANSPORT NOT a_LC6_E16  ;
and2_3328: n_3979 <=  n_3980  AND n_3981;
delay_3329: n_3980  <= TRANSPORT a_N965  ;
delay_3330: n_3981  <= TRANSPORT a_LC6_E5  ;
and1_3331: n_3982 <=  gnd;
dff_3332: DFF_a8237

    PORT MAP ( D => a_EQ1155, CLK => a_SH3WRDCNTREG_F14_G_aCLK, CLRN => a_SH3WRDCNTREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SH3WRDCNTREG_F14_G);
inv_3333: a_SH3WRDCNTREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3334: a_EQ1155 <=  n_3989  XOR n_3996;
or2_3335: n_3989 <=  n_3990  OR n_3993;
and2_3336: n_3990 <=  n_3991  AND n_3992;
inv_3337: n_3991  <= TRANSPORT NOT a_N2528  ;
delay_3338: n_3992  <= TRANSPORT a_LC5_E5  ;
and2_3339: n_3993 <=  n_3994  AND n_3995;
delay_3340: n_3994  <= TRANSPORT a_SCH3BWORDOUT_F14_G  ;
delay_3341: n_3995  <= TRANSPORT a_N2528  ;
and1_3342: n_3996 <=  gnd;
delay_3343: n_3997  <= TRANSPORT clk  ;
filter_3344: FILTER_a8237

    PORT MAP (IN1 => n_3997, Y => a_SH3WRDCNTREG_F14_G_aCLK);
delay_3345: a_N869_aNOT  <= TRANSPORT a_EQ318  ;
xor2_3346: a_EQ318 <=  n_4001  XOR n_4009;
or2_3347: n_4001 <=  n_4002  OR n_4005;
and2_3348: n_4002 <=  n_4003  AND n_4004;
inv_3349: n_4003  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_3350: n_4004  <= TRANSPORT dbin(6)  ;
and2_3351: n_4005 <=  n_4006  AND n_4007;
delay_3352: n_4006  <= TRANSPORT a_N2577_aNOT  ;
delay_3353: n_4007  <= TRANSPORT a_SH1WRDCNTREG_F14_G  ;
and1_3354: n_4009 <=  gnd;
delay_3355: a_LC7_E19  <= TRANSPORT a_EQ316  ;
xor2_3356: a_EQ316 <=  n_4012  XOR n_4019;
or2_3357: n_4012 <=  n_4013  OR n_4016;
and2_3358: n_4013 <=  n_4014  AND n_4015;
inv_3359: n_4014  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_3360: n_4015  <= TRANSPORT NOT a_LC6_E16  ;
and2_3361: n_4016 <=  n_4017  AND n_4018;
delay_3362: n_4017  <= TRANSPORT a_N2559_aNOT  ;
delay_3363: n_4018  <= TRANSPORT a_N869_aNOT  ;
and1_3364: n_4019 <=  gnd;
dff_3365: DFF_a8237

    PORT MAP ( D => a_EQ1143, CLK => a_SH1WRDCNTREG_F14_G_aCLK, CLRN => a_SH1WRDCNTREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SH1WRDCNTREG_F14_G);
inv_3366: a_SH1WRDCNTREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3367: a_EQ1143 <=  n_4026  XOR n_4033;
or2_3368: n_4026 <=  n_4027  OR n_4030;
and2_3369: n_4027 <=  n_4028  AND n_4029;
delay_3370: n_4028  <= TRANSPORT a_SCH1BWORDOUT_F14_G  ;
delay_3371: n_4029  <= TRANSPORT a_N2526  ;
and2_3372: n_4030 <=  n_4031  AND n_4032;
inv_3373: n_4031  <= TRANSPORT NOT a_N2526  ;
delay_3374: n_4032  <= TRANSPORT a_LC7_E19  ;
and1_3375: n_4033 <=  gnd;
delay_3376: n_4034  <= TRANSPORT clk  ;
filter_3377: FILTER_a8237

    PORT MAP (IN1 => n_4034, Y => a_SH1WRDCNTREG_F14_G_aCLK);
delay_3378: a_LC8_E4  <= TRANSPORT a_EQ314  ;
xor2_3379: a_EQ314 <=  n_4038  XOR n_4050;
or3_3380: n_4038 <=  n_4039  OR n_4043  OR n_4047;
and3_3381: n_4039 <=  n_4040  AND n_4041  AND n_4042;
inv_3382: n_4040  <= TRANSPORT NOT a_LC3_D22  ;
inv_3383: n_4041  <= TRANSPORT NOT a_N62_aNOT  ;
delay_3384: n_4042  <= TRANSPORT dbin(6)  ;
and2_3385: n_4043 <=  n_4044  AND n_4045;
delay_3386: n_4044  <= TRANSPORT a_N62_aNOT  ;
delay_3387: n_4045  <= TRANSPORT a_SH2WRDCNTREG_F14_G  ;
and2_3388: n_4047 <=  n_4048  AND n_4049;
delay_3389: n_4048  <= TRANSPORT a_LC3_D22  ;
delay_3390: n_4049  <= TRANSPORT a_SH2WRDCNTREG_F14_G  ;
and1_3391: n_4050 <=  gnd;
delay_3392: a_LC7_E4  <= TRANSPORT a_EQ323  ;
xor2_3393: a_EQ323 <=  n_4053  XOR n_4060;
or2_3394: n_4053 <=  n_4054  OR n_4057;
and2_3395: n_4054 <=  n_4055  AND n_4056;
inv_3396: n_4055  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_3397: n_4056  <= TRANSPORT NOT a_LC6_E16  ;
and2_3398: n_4057 <=  n_4058  AND n_4059;
delay_3399: n_4058  <= TRANSPORT a_N2560_aNOT  ;
delay_3400: n_4059  <= TRANSPORT a_LC8_E4  ;
and1_3401: n_4060 <=  gnd;
dff_3402: DFF_a8237

    PORT MAP ( D => a_EQ1149, CLK => a_SH2WRDCNTREG_F14_G_aCLK, CLRN => a_SH2WRDCNTREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SH2WRDCNTREG_F14_G);
inv_3403: a_SH2WRDCNTREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3404: a_EQ1149 <=  n_4067  XOR n_4074;
or2_3405: n_4067 <=  n_4068  OR n_4071;
and2_3406: n_4068 <=  n_4069  AND n_4070;
inv_3407: n_4069  <= TRANSPORT NOT a_N2527  ;
delay_3408: n_4070  <= TRANSPORT a_LC7_E4  ;
and2_3409: n_4071 <=  n_4072  AND n_4073;
delay_3410: n_4072  <= TRANSPORT a_SCH2BWORDOUT_F14_G  ;
delay_3411: n_4073  <= TRANSPORT a_N2527  ;
and1_3412: n_4074 <=  gnd;
delay_3413: n_4075  <= TRANSPORT clk  ;
filter_3414: FILTER_a8237

    PORT MAP (IN1 => n_4075, Y => a_SH2WRDCNTREG_F14_G_aCLK);
delay_3415: a_LC2_E13  <= TRANSPORT a_EQ750  ;
xor2_3416: a_EQ750 <=  n_4079  XOR n_4091;
or3_3417: n_4079 <=  n_4080  OR n_4084  OR n_4088;
and3_3418: n_4080 <=  n_4081  AND n_4082  AND n_4083;
inv_3419: n_4081  <= TRANSPORT NOT a_LC3_D22  ;
inv_3420: n_4082  <= TRANSPORT NOT a_N2353  ;
delay_3421: n_4083  <= TRANSPORT dbin(6)  ;
and2_3422: n_4084 <=  n_4085  AND n_4086;
delay_3423: n_4085  <= TRANSPORT a_N2353  ;
delay_3424: n_4086  <= TRANSPORT a_SH0WRDCNTREG_F14_G  ;
and2_3425: n_4088 <=  n_4089  AND n_4090;
delay_3426: n_4089  <= TRANSPORT a_LC3_D22  ;
delay_3427: n_4090  <= TRANSPORT a_SH0WRDCNTREG_F14_G  ;
and1_3428: n_4091 <=  gnd;
delay_3429: a_LC3_E13  <= TRANSPORT a_EQ751  ;
xor2_3430: a_EQ751 <=  n_4094  XOR n_4101;
or2_3431: n_4094 <=  n_4095  OR n_4098;
and2_3432: n_4095 <=  n_4096  AND n_4097;
inv_3433: n_4096  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_3434: n_4097  <= TRANSPORT NOT a_LC6_E16  ;
and2_3435: n_4098 <=  n_4099  AND n_4100;
delay_3436: n_4099  <= TRANSPORT a_N2558_aNOT  ;
delay_3437: n_4100  <= TRANSPORT a_LC2_E13  ;
and1_3438: n_4101 <=  gnd;
dff_3439: DFF_a8237

    PORT MAP ( D => a_EQ1137, CLK => a_SH0WRDCNTREG_F14_G_aCLK, CLRN => a_SH0WRDCNTREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SH0WRDCNTREG_F14_G);
inv_3440: a_SH0WRDCNTREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3441: a_EQ1137 <=  n_4108  XOR n_4115;
or2_3442: n_4108 <=  n_4109  OR n_4112;
and2_3443: n_4109 <=  n_4110  AND n_4111;
inv_3444: n_4110  <= TRANSPORT NOT a_N2525  ;
delay_3445: n_4111  <= TRANSPORT a_LC3_E13  ;
and2_3446: n_4112 <=  n_4113  AND n_4114;
delay_3447: n_4113  <= TRANSPORT a_SCH0BWORDOUT_F14_G  ;
delay_3448: n_4114  <= TRANSPORT a_N2525  ;
and1_3449: n_4115 <=  gnd;
delay_3450: n_4116  <= TRANSPORT clk  ;
filter_3451: FILTER_a8237

    PORT MAP (IN1 => n_4116, Y => a_SH0WRDCNTREG_F14_G_aCLK);
delay_3452: a_LC2_C25  <= TRANSPORT a_EQ399  ;
xor2_3453: a_EQ399 <=  n_4120  XOR n_4127;
or2_3454: n_4120 <=  n_4121  OR n_4124;
and2_3455: n_4121 <=  n_4122  AND n_4123;
inv_3456: n_4122  <= TRANSPORT NOT a_N88_aNOT  ;
delay_3457: n_4123  <= TRANSPORT a_SCH1WRDCNTREG_F4_G  ;
and2_3458: n_4124 <=  n_4125  AND n_4126;
inv_3459: n_4125  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_3460: n_4126  <= TRANSPORT a_SCH0WRDCNTREG_F4_G  ;
and1_3461: n_4127 <=  gnd;
delay_3462: a_N1296_aNOT  <= TRANSPORT a_EQ409  ;
xor2_3463: a_EQ409 <=  n_4130  XOR n_4141;
or3_3464: n_4130 <=  n_4131  OR n_4135  OR n_4138;
and3_3465: n_4131 <=  n_4132  AND n_4133  AND n_4134;
delay_3466: n_4132  <= TRANSPORT a_N2557  ;
inv_3467: n_4133  <= TRANSPORT NOT a_LC3_C13  ;
inv_3468: n_4134  <= TRANSPORT NOT a_N3552  ;
and2_3469: n_4135 <=  n_4136  AND n_4137;
delay_3470: n_4136  <= TRANSPORT a_LC3_C13  ;
delay_3471: n_4137  <= TRANSPORT a_N3552  ;
and2_3472: n_4138 <=  n_4139  AND n_4140;
inv_3473: n_4139  <= TRANSPORT NOT a_N2557  ;
delay_3474: n_4140  <= TRANSPORT a_N3552  ;
and1_3475: n_4141 <=  gnd;
delay_3476: a_N1280  <= TRANSPORT a_EQ398  ;
xor2_3477: a_EQ398 <=  n_4144  XOR n_4151;
or2_3478: n_4144 <=  n_4145  OR n_4148;
and2_3479: n_4145 <=  n_4146  AND n_4147;
delay_3480: n_4146  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_3481: n_4147  <= TRANSPORT a_SCH1WRDCNTREG_F4_G  ;
and2_3482: n_4148 <=  n_4149  AND n_4150;
inv_3483: n_4149  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_3484: n_4150  <= TRANSPORT a_SCH0WRDCNTREG_F4_G  ;
and1_3485: n_4151 <=  gnd;
delay_3486: a_N1279  <= TRANSPORT a_EQ397  ;
xor2_3487: a_EQ397 <=  n_4154  XOR n_4163;
or3_3488: n_4154 <=  n_4155  OR n_4157  OR n_4160;
and1_3489: n_4155 <=  n_4156;
delay_3490: n_4156  <= TRANSPORT startdma  ;
and2_3491: n_4157 <=  n_4158  AND n_4159;
inv_3492: n_4158  <= TRANSPORT NOT a_N2531  ;
delay_3493: n_4159  <= TRANSPORT a_N1296_aNOT  ;
and2_3494: n_4160 <=  n_4161  AND n_4162;
delay_3495: n_4161  <= TRANSPORT a_N2531  ;
delay_3496: n_4162  <= TRANSPORT a_N1280  ;
and1_3497: n_4163 <=  gnd;
delay_3498: a_LC3_C25  <= TRANSPORT a_EQ400  ;
xor2_3499: a_EQ400 <=  n_4166  XOR n_4173;
or2_3500: n_4166 <=  n_4167  OR n_4170;
and2_3501: n_4167 <=  n_4168  AND n_4169;
inv_3502: n_4168  <= TRANSPORT NOT a_N2376  ;
delay_3503: n_4169  <= TRANSPORT a_SCH2WRDCNTREG_F4_G  ;
and2_3504: n_4170 <=  n_4171  AND n_4172;
inv_3505: n_4171  <= TRANSPORT NOT a_N2377  ;
delay_3506: n_4172  <= TRANSPORT a_SCH3WRDCNTREG_F4_G  ;
and1_3507: n_4173 <=  gnd;
dff_3508: DFF_a8237

    PORT MAP ( D => a_EQ848, CLK => a_N3552_aCLK, CLRN => a_N3552_aCLRN, PRN => vcc,
          Q => a_N3552);
inv_3509: a_N3552_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3510: a_EQ848 <=  n_4180  XOR n_4190;
or3_3511: n_4180 <=  n_4181  OR n_4184  OR n_4187;
and2_3512: n_4181 <=  n_4182  AND n_4183;
delay_3513: n_4182  <= TRANSPORT a_LC2_C25  ;
delay_3514: n_4183  <= TRANSPORT a_N1279  ;
and2_3515: n_4184 <=  n_4185  AND n_4186;
delay_3516: n_4185  <= TRANSPORT a_N1279  ;
inv_3517: n_4186  <= TRANSPORT NOT startdma  ;
and2_3518: n_4187 <=  n_4188  AND n_4189;
delay_3519: n_4188  <= TRANSPORT a_N1279  ;
delay_3520: n_4189  <= TRANSPORT a_LC3_C25  ;
and1_3521: n_4190 <=  gnd;
delay_3522: n_4191  <= TRANSPORT clk  ;
filter_3523: FILTER_a8237

    PORT MAP (IN1 => n_4191, Y => a_N3552_aCLK);
delay_3524: a_LC6_F16  <= TRANSPORT a_EQ268  ;
xor2_3525: a_EQ268 <=  n_4195  XOR n_4210;
or4_3526: n_4195 <=  n_4196  OR n_4199  OR n_4202  OR n_4205;
and2_3527: n_4196 <=  n_4197  AND n_4198;
delay_3528: n_4197  <= TRANSPORT a_N3552  ;
delay_3529: n_4198  <= TRANSPORT a_N3551  ;
and2_3530: n_4199 <=  n_4200  AND n_4201;
delay_3531: n_4200  <= TRANSPORT a_LC3_C13  ;
delay_3532: n_4201  <= TRANSPORT a_N3551  ;
and2_3533: n_4202 <=  n_4203  AND n_4204;
inv_3534: n_4203  <= TRANSPORT NOT a_N2557  ;
delay_3535: n_4204  <= TRANSPORT a_N3551  ;
and4_3536: n_4205 <=  n_4206  AND n_4207  AND n_4208  AND n_4209;
delay_3537: n_4206  <= TRANSPORT a_N2557  ;
inv_3538: n_4207  <= TRANSPORT NOT a_LC3_C13  ;
inv_3539: n_4208  <= TRANSPORT NOT a_N3552  ;
inv_3540: n_4209  <= TRANSPORT NOT a_N3551  ;
and1_3541: n_4210 <=  gnd;
delay_3542: a_LC4_F16  <= TRANSPORT a_EQ267  ;
xor2_3543: a_EQ267 <=  n_4213  XOR n_4222;
or2_3544: n_4213 <=  n_4214  OR n_4218;
and2_3545: n_4214 <=  n_4215  AND n_4216;
delay_3546: n_4215  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_3547: n_4216  <= TRANSPORT a_SCH1WRDCNTREG_F5_G  ;
and2_3548: n_4218 <=  n_4219  AND n_4220;
inv_3549: n_4219  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_3550: n_4220  <= TRANSPORT a_SCH0WRDCNTREG_F5_G  ;
and1_3551: n_4222 <=  gnd;
delay_3552: a_N522_aNOT  <= TRANSPORT a_EQ264  ;
xor2_3553: a_EQ264 <=  n_4225  XOR n_4232;
or2_3554: n_4225 <=  n_4226  OR n_4229;
and2_3555: n_4226 <=  n_4227  AND n_4228;
inv_3556: n_4227  <= TRANSPORT NOT a_N2531  ;
delay_3557: n_4228  <= TRANSPORT a_LC6_F16  ;
and2_3558: n_4229 <=  n_4230  AND n_4231;
delay_3559: n_4230  <= TRANSPORT a_N2531  ;
delay_3560: n_4231  <= TRANSPORT a_LC4_F16  ;
and1_3561: n_4232 <=  gnd;
delay_3562: a_LC3_F16  <= TRANSPORT a_EQ266  ;
xor2_3563: a_EQ266 <=  n_4235  XOR n_4243;
or2_3564: n_4235 <=  n_4236  OR n_4240;
and2_3565: n_4236 <=  n_4237  AND n_4238;
inv_3566: n_4237  <= TRANSPORT NOT a_N2376  ;
delay_3567: n_4238  <= TRANSPORT a_SCH2WRDCNTREG_F5_G  ;
and2_3568: n_4240 <=  n_4241  AND n_4242;
inv_3569: n_4241  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_3570: n_4242  <= TRANSPORT a_SCH0WRDCNTREG_F5_G  ;
and1_3571: n_4243 <=  gnd;
delay_3572: a_LC1_F16  <= TRANSPORT a_EQ265  ;
xor2_3573: a_EQ265 <=  n_4246  XOR n_4254;
or2_3574: n_4246 <=  n_4247  OR n_4250;
and2_3575: n_4247 <=  n_4248  AND n_4249;
inv_3576: n_4248  <= TRANSPORT NOT a_N88_aNOT  ;
delay_3577: n_4249  <= TRANSPORT a_SCH1WRDCNTREG_F5_G  ;
and2_3578: n_4250 <=  n_4251  AND n_4252;
inv_3579: n_4251  <= TRANSPORT NOT a_N2377  ;
delay_3580: n_4252  <= TRANSPORT a_SCH3WRDCNTREG_F5_G  ;
and1_3581: n_4254 <=  gnd;
dff_3582: DFF_a8237

    PORT MAP ( D => a_EQ847, CLK => a_N3551_aCLK, CLRN => a_N3551_aCLRN, PRN => vcc,
          Q => a_N3551);
inv_3583: a_N3551_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3584: a_EQ847 <=  n_4261  XOR n_4271;
or3_3585: n_4261 <=  n_4262  OR n_4265  OR n_4268;
and2_3586: n_4262 <=  n_4263  AND n_4264;
delay_3587: n_4263  <= TRANSPORT a_N522_aNOT  ;
inv_3588: n_4264  <= TRANSPORT NOT startdma  ;
and2_3589: n_4265 <=  n_4266  AND n_4267;
delay_3590: n_4266  <= TRANSPORT a_LC3_F16  ;
delay_3591: n_4267  <= TRANSPORT startdma  ;
and2_3592: n_4268 <=  n_4269  AND n_4270;
delay_3593: n_4269  <= TRANSPORT a_LC1_F16  ;
delay_3594: n_4270  <= TRANSPORT startdma  ;
and1_3595: n_4271 <=  gnd;
delay_3596: n_4272  <= TRANSPORT clk  ;
filter_3597: FILTER_a8237

    PORT MAP (IN1 => n_4272, Y => a_N3551_aCLK);
delay_3598: a_LC6_F13  <= TRANSPORT a_EQ505  ;
xor2_3599: a_EQ505 <=  n_4276  XOR n_4283;
or2_3600: n_4276 <=  n_4277  OR n_4280;
and2_3601: n_4277 <=  n_4278  AND n_4279;
inv_3602: n_4278  <= TRANSPORT NOT a_N2557  ;
delay_3603: n_4279  <= TRANSPORT a_N3550  ;
and2_3604: n_4280 <=  n_4281  AND n_4282;
delay_3605: n_4281  <= TRANSPORT a_N2557  ;
inv_3606: n_4282  <= TRANSPORT NOT a_LC7_F13  ;
and1_3607: n_4283 <=  gnd;
delay_3608: a_LC5_F13  <= TRANSPORT a_EQ504  ;
xor2_3609: a_EQ504 <=  n_4286  XOR n_4293;
or2_3610: n_4286 <=  n_4287  OR n_4290;
and2_3611: n_4287 <=  n_4288  AND n_4289;
inv_3612: n_4288  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_3613: n_4289  <= TRANSPORT a_SCH0WRDCNTREG_F6_G  ;
and2_3614: n_4290 <=  n_4291  AND n_4292;
delay_3615: n_4291  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_3616: n_4292  <= TRANSPORT a_SCH1WRDCNTREG_F6_G  ;
and1_3617: n_4293 <=  gnd;
delay_3618: a_N1764_aNOT  <= TRANSPORT a_EQ506  ;
xor2_3619: a_EQ506 <=  n_4296  XOR n_4303;
or2_3620: n_4296 <=  n_4297  OR n_4300;
and2_3621: n_4297 <=  n_4298  AND n_4299;
inv_3622: n_4298  <= TRANSPORT NOT a_N2531  ;
delay_3623: n_4299  <= TRANSPORT a_LC6_F13  ;
and2_3624: n_4300 <=  n_4301  AND n_4302;
delay_3625: n_4301  <= TRANSPORT a_N2531  ;
delay_3626: n_4302  <= TRANSPORT a_LC5_F13  ;
and1_3627: n_4303 <=  gnd;
delay_3628: a_LC1_F13  <= TRANSPORT a_EQ503  ;
xor2_3629: a_EQ503 <=  n_4306  XOR n_4313;
or2_3630: n_4306 <=  n_4307  OR n_4310;
and2_3631: n_4307 <=  n_4308  AND n_4309;
inv_3632: n_4308  <= TRANSPORT NOT a_N88_aNOT  ;
delay_3633: n_4309  <= TRANSPORT a_SCH1WRDCNTREG_F6_G  ;
and2_3634: n_4310 <=  n_4311  AND n_4312;
inv_3635: n_4311  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_3636: n_4312  <= TRANSPORT a_SCH0WRDCNTREG_F6_G  ;
and1_3637: n_4313 <=  gnd;
delay_3638: a_LC2_F13  <= TRANSPORT a_EQ502  ;
xor2_3639: a_EQ502 <=  n_4316  XOR n_4323;
or2_3640: n_4316 <=  n_4317  OR n_4320;
and2_3641: n_4317 <=  n_4318  AND n_4319;
inv_3642: n_4318  <= TRANSPORT NOT a_N2376  ;
delay_3643: n_4319  <= TRANSPORT a_SCH2WRDCNTREG_F6_G  ;
and2_3644: n_4320 <=  n_4321  AND n_4322;
inv_3645: n_4321  <= TRANSPORT NOT a_N2377  ;
delay_3646: n_4322  <= TRANSPORT a_SCH3WRDCNTREG_F6_G  ;
and1_3647: n_4323 <=  gnd;
dff_3648: DFF_a8237

    PORT MAP ( D => a_EQ846, CLK => a_N3550_aCLK, CLRN => a_N3550_aCLRN, PRN => vcc,
          Q => a_N3550);
inv_3649: a_N3550_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3650: a_EQ846 <=  n_4330  XOR n_4340;
or3_3651: n_4330 <=  n_4331  OR n_4334  OR n_4337;
and2_3652: n_4331 <=  n_4332  AND n_4333;
delay_3653: n_4332  <= TRANSPORT a_N1764_aNOT  ;
inv_3654: n_4333  <= TRANSPORT NOT startdma  ;
and2_3655: n_4334 <=  n_4335  AND n_4336;
delay_3656: n_4335  <= TRANSPORT a_LC1_F13  ;
delay_3657: n_4336  <= TRANSPORT startdma  ;
and2_3658: n_4337 <=  n_4338  AND n_4339;
delay_3659: n_4338  <= TRANSPORT a_LC2_F13  ;
delay_3660: n_4339  <= TRANSPORT startdma  ;
and1_3661: n_4340 <=  gnd;
delay_3662: n_4341  <= TRANSPORT clk  ;
filter_3663: FILTER_a8237

    PORT MAP (IN1 => n_4341, Y => a_N3550_aCLK);
delay_3664: a_LC1_E11  <= TRANSPORT a_EQ518  ;
xor2_3665: a_EQ518 <=  n_4345  XOR n_4354;
or2_3666: n_4345 <=  n_4346  OR n_4350;
and2_3667: n_4346 <=  n_4347  AND n_4348;
inv_3668: n_4347  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_3669: n_4348  <= TRANSPORT a_SCH0MODEREG_F3_G  ;
and2_3670: n_4350 <=  n_4351  AND n_4352;
inv_3671: n_4351  <= TRANSPORT NOT a_N88_aNOT  ;
delay_3672: n_4352  <= TRANSPORT a_SCH1MODEREG_F3_G  ;
and1_3673: n_4354 <=  gnd;
delay_3674: a_N1879_aNOT  <= TRANSPORT a_EQ517  ;
xor2_3675: a_EQ517 <=  n_4357  XOR n_4366;
or3_3676: n_4357 <=  n_4358  OR n_4361  OR n_4364;
and2_3677: n_4358 <=  n_4359  AND n_4360;
delay_3678: n_4359  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_3679: n_4360  <= TRANSPORT a_SCH0MODEREG_F3_G  ;
and2_3680: n_4361 <=  n_4362  AND n_4363;
inv_3681: n_4362  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_3682: n_4363  <= TRANSPORT a_SCH1MODEREG_F3_G  ;
and1_3683: n_4364 <=  n_4365;
inv_3684: n_4365  <= TRANSPORT NOT a_N2591  ;
and1_3685: n_4366 <=  gnd;
delay_3686: a_LC1_E1  <= TRANSPORT a_EQ589  ;
xor2_3687: a_EQ589 <=  n_4369  XOR n_4378;
or2_3688: n_4369 <=  n_4370  OR n_4374;
and2_3689: n_4370 <=  n_4371  AND n_4372;
inv_3690: n_4371  <= TRANSPORT NOT a_N2377  ;
delay_3691: n_4372  <= TRANSPORT a_SCH3MODEREG_F3_G  ;
and2_3692: n_4374 <=  n_4375  AND n_4376;
inv_3693: n_4375  <= TRANSPORT NOT a_N2376  ;
delay_3694: n_4376  <= TRANSPORT a_SCH2MODEREG_F3_G  ;
and1_3695: n_4378 <=  gnd;
delay_3696: a_N2529  <= TRANSPORT a_EQ590  ;
xor2_3697: a_EQ590 <=  n_4381  XOR n_4390;
or3_3698: n_4381 <=  n_4382  OR n_4385  OR n_4388;
and2_3699: n_4382 <=  n_4383  AND n_4384;
delay_3700: n_4383  <= TRANSPORT a_LC1_E11  ;
delay_3701: n_4384  <= TRANSPORT a_N1879_aNOT  ;
and2_3702: n_4385 <=  n_4386  AND n_4387;
delay_3703: n_4386  <= TRANSPORT a_N2591  ;
delay_3704: n_4387  <= TRANSPORT a_N1879_aNOT  ;
and1_3705: n_4388 <=  n_4389;
delay_3706: n_4389  <= TRANSPORT a_LC1_E1  ;
and1_3707: n_4390 <=  gnd;
delay_3708: a_N2530_aNOT  <= TRANSPORT a_EQ591  ;
xor2_3709: a_EQ591 <=  n_4393  XOR n_4399;
or2_3710: n_4393 <=  n_4394  OR n_4397;
and1_3711: n_4394 <=  n_4395;
inv_3712: n_4395  <= TRANSPORT NOT a_SCOMMANDREG_F1_G  ;
and1_3713: n_4397 <=  n_4398;
delay_3714: n_4398  <= TRANSPORT a_N2598_aNOT  ;
and1_3715: n_4399 <=  gnd;
delay_3716: a_N757  <= TRANSPORT a_N757_aIN  ;
xor2_3717: a_N757_aIN <=  n_4402  XOR n_4406;
or1_3718: n_4402 <=  n_4403;
and2_3719: n_4403 <=  n_4404  AND n_4405;
delay_3720: n_4404  <= TRANSPORT a_N2529  ;
delay_3721: n_4405  <= TRANSPORT a_N2530_aNOT  ;
and1_3722: n_4406 <=  gnd;
delay_3723: a_LC2_C14  <= TRANSPORT a_EQ002  ;
xor2_3724: a_EQ002 <=  n_4409  XOR n_4434;
or6_3725: n_4409 <=  n_4410  OR n_4414  OR n_4418  OR n_4422  OR n_4426  OR n_4430;
and3_3726: n_4410 <=  n_4411  AND n_4412  AND n_4413;
delay_3727: n_4411  <= TRANSPORT a_LC7_D18  ;
delay_3728: n_4412  <= TRANSPORT a_LC7_C17  ;
inv_3729: n_4413  <= TRANSPORT NOT a_LC4_C16  ;
and3_3730: n_4414 <=  n_4415  AND n_4416  AND n_4417;
delay_3731: n_4415  <= TRANSPORT a_N757  ;
delay_3732: n_4416  <= TRANSPORT a_LC7_D18  ;
inv_3733: n_4417  <= TRANSPORT NOT a_LC4_C16  ;
and3_3734: n_4418 <=  n_4419  AND n_4420  AND n_4421;
delay_3735: n_4419  <= TRANSPORT a_N757  ;
delay_3736: n_4420  <= TRANSPORT a_LC7_C17  ;
inv_3737: n_4421  <= TRANSPORT NOT a_LC4_C16  ;
and3_3738: n_4422 <=  n_4423  AND n_4424  AND n_4425;
inv_3739: n_4423  <= TRANSPORT NOT a_N757  ;
inv_3740: n_4424  <= TRANSPORT NOT a_LC7_C17  ;
delay_3741: n_4425  <= TRANSPORT a_LC4_C16  ;
and3_3742: n_4426 <=  n_4427  AND n_4428  AND n_4429;
inv_3743: n_4427  <= TRANSPORT NOT a_N757  ;
inv_3744: n_4428  <= TRANSPORT NOT a_LC7_D18  ;
delay_3745: n_4429  <= TRANSPORT a_LC4_C16  ;
and3_3746: n_4430 <=  n_4431  AND n_4432  AND n_4433;
inv_3747: n_4431  <= TRANSPORT NOT a_LC7_D18  ;
inv_3748: n_4432  <= TRANSPORT NOT a_LC7_C17  ;
delay_3749: n_4433  <= TRANSPORT a_LC4_C16  ;
and1_3750: n_4434 <=  gnd;
delay_3751: a_LC6_C14  <= TRANSPORT a_LC6_C14_aIN  ;
xor2_3752: a_LC6_C14_aIN <=  n_4437  XOR n_4447;
or3_3753: n_4437 <=  n_4438  OR n_4441  OR n_4444;
and2_3754: n_4438 <=  n_4439  AND n_4440;
delay_3755: n_4439  <= TRANSPORT a_LC7_D18  ;
delay_3756: n_4440  <= TRANSPORT a_LC7_C17  ;
and2_3757: n_4441 <=  n_4442  AND n_4443;
delay_3758: n_4442  <= TRANSPORT a_N757  ;
delay_3759: n_4443  <= TRANSPORT a_LC7_D18  ;
and2_3760: n_4444 <=  n_4445  AND n_4446;
delay_3761: n_4445  <= TRANSPORT a_N757  ;
delay_3762: n_4446  <= TRANSPORT a_LC7_C17  ;
and1_3763: n_4447 <=  gnd;
delay_3764: a_LC3_C14  <= TRANSPORT a_EQ019  ;
xor2_3765: a_EQ019 <=  n_4450  XOR n_4457;
or2_3766: n_4450 <=  n_4451  OR n_4454;
and2_3767: n_4451 <=  n_4452  AND n_4453;
delay_3768: n_4452  <= TRANSPORT a_N757  ;
delay_3769: n_4453  <= TRANSPORT a_LC2_C14  ;
and2_3770: n_4454 <=  n_4455  AND n_4456;
delay_3771: n_4455  <= TRANSPORT a_LC6_C14  ;
delay_3772: n_4456  <= TRANSPORT a_LC4_C16  ;
and1_3773: n_4457 <=  gnd;
delay_3774: a_LC4_C14  <= TRANSPORT a_EQ021  ;
xor2_3775: a_EQ021 <=  n_4460  XOR n_4474;
or4_3776: n_4460 <=  n_4461  OR n_4464  OR n_4467  OR n_4470;
and2_3777: n_4461 <=  n_4462  AND n_4463;
delay_3778: n_4462  <= TRANSPORT a_N757  ;
delay_3779: n_4463  <= TRANSPORT a_LC4_C16  ;
and2_3780: n_4464 <=  n_4465  AND n_4466;
delay_3781: n_4465  <= TRANSPORT a_N757  ;
delay_3782: n_4466  <= TRANSPORT a_LC7_C17  ;
and2_3783: n_4467 <=  n_4468  AND n_4469;
delay_3784: n_4468  <= TRANSPORT a_N757  ;
delay_3785: n_4469  <= TRANSPORT a_LC7_D18  ;
and3_3786: n_4470 <=  n_4471  AND n_4472  AND n_4473;
delay_3787: n_4471  <= TRANSPORT a_LC7_D18  ;
delay_3788: n_4472  <= TRANSPORT a_LC7_C17  ;
delay_3789: n_4473  <= TRANSPORT a_LC4_C16  ;
and1_3790: n_4474 <=  gnd;
delay_3791: a_LC7_C14  <= TRANSPORT a_EQ020  ;
xor2_3792: a_EQ020 <=  n_4477  XOR n_4489;
or3_3793: n_4477 <=  n_4478  OR n_4481  OR n_4485;
and2_3794: n_4478 <=  n_4479  AND n_4480;
delay_3795: n_4479  <= TRANSPORT a_LC3_C14  ;
delay_3796: n_4480  <= TRANSPORT a_LC2_C24  ;
and3_3797: n_4481 <=  n_4482  AND n_4483  AND n_4484;
delay_3798: n_4482  <= TRANSPORT a_N757  ;
inv_3799: n_4483  <= TRANSPORT NOT a_LC4_C14  ;
delay_3800: n_4484  <= TRANSPORT a_LC2_C24  ;
and3_3801: n_4485 <=  n_4486  AND n_4487  AND n_4488;
delay_3802: n_4486  <= TRANSPORT a_N757  ;
delay_3803: n_4487  <= TRANSPORT a_LC4_C14  ;
inv_3804: n_4488  <= TRANSPORT NOT a_LC2_C24  ;
and1_3805: n_4489 <=  gnd;
delay_3806: a_LC1_F26  <= TRANSPORT a_EQ003  ;
xor2_3807: a_EQ003 <=  n_4492  XOR n_4517;
or6_3808: n_4492 <=  n_4493  OR n_4497  OR n_4501  OR n_4505  OR n_4509  OR n_4513;
and3_3809: n_4493 <=  n_4494  AND n_4495  AND n_4496;
delay_3810: n_4494  <= TRANSPORT a_LC7_C14  ;
delay_3811: n_4495  <= TRANSPORT a_LC1_C16  ;
inv_3812: n_4496  <= TRANSPORT NOT a_LC3_F6  ;
and3_3813: n_4497 <=  n_4498  AND n_4499  AND n_4500;
delay_3814: n_4498  <= TRANSPORT a_N757  ;
delay_3815: n_4499  <= TRANSPORT a_LC7_C14  ;
inv_3816: n_4500  <= TRANSPORT NOT a_LC3_F6  ;
and3_3817: n_4501 <=  n_4502  AND n_4503  AND n_4504;
delay_3818: n_4502  <= TRANSPORT a_N757  ;
delay_3819: n_4503  <= TRANSPORT a_LC1_C16  ;
inv_3820: n_4504  <= TRANSPORT NOT a_LC3_F6  ;
and3_3821: n_4505 <=  n_4506  AND n_4507  AND n_4508;
inv_3822: n_4506  <= TRANSPORT NOT a_N757  ;
inv_3823: n_4507  <= TRANSPORT NOT a_LC1_C16  ;
delay_3824: n_4508  <= TRANSPORT a_LC3_F6  ;
and3_3825: n_4509 <=  n_4510  AND n_4511  AND n_4512;
inv_3826: n_4510  <= TRANSPORT NOT a_N757  ;
inv_3827: n_4511  <= TRANSPORT NOT a_LC7_C14  ;
delay_3828: n_4512  <= TRANSPORT a_LC3_F6  ;
and3_3829: n_4513 <=  n_4514  AND n_4515  AND n_4516;
inv_3830: n_4514  <= TRANSPORT NOT a_LC7_C14  ;
inv_3831: n_4515  <= TRANSPORT NOT a_LC1_C16  ;
delay_3832: n_4516  <= TRANSPORT a_LC3_F6  ;
and1_3833: n_4517 <=  gnd;
delay_3834: a_LC4_F20  <= TRANSPORT a_LC4_F20_aIN  ;
xor2_3835: a_LC4_F20_aIN <=  n_4520  XOR n_4530;
or3_3836: n_4520 <=  n_4521  OR n_4524  OR n_4527;
and2_3837: n_4521 <=  n_4522  AND n_4523;
delay_3838: n_4522  <= TRANSPORT a_LC7_C14  ;
delay_3839: n_4523  <= TRANSPORT a_LC1_C16  ;
and2_3840: n_4524 <=  n_4525  AND n_4526;
delay_3841: n_4525  <= TRANSPORT a_N757  ;
delay_3842: n_4526  <= TRANSPORT a_LC7_C14  ;
and2_3843: n_4527 <=  n_4528  AND n_4529;
delay_3844: n_4528  <= TRANSPORT a_N757  ;
delay_3845: n_4529  <= TRANSPORT a_LC1_C16  ;
and1_3846: n_4530 <=  gnd;
delay_3847: a_LC6_F20  <= TRANSPORT a_EQ017  ;
xor2_3848: a_EQ017 <=  n_4533  XOR n_4540;
or2_3849: n_4533 <=  n_4534  OR n_4537;
and2_3850: n_4534 <=  n_4535  AND n_4536;
delay_3851: n_4535  <= TRANSPORT a_N757  ;
delay_3852: n_4536  <= TRANSPORT a_LC1_F26  ;
and2_3853: n_4537 <=  n_4538  AND n_4539;
delay_3854: n_4538  <= TRANSPORT a_LC4_F20  ;
delay_3855: n_4539  <= TRANSPORT a_LC3_F6  ;
and1_3856: n_4540 <=  gnd;
delay_3857: a_LC6_F15  <= TRANSPORT a_EQ016  ;
xor2_3858: a_EQ016 <=  n_4543  XOR n_4553;
or3_3859: n_4543 <=  n_4544  OR n_4547  OR n_4550;
and2_3860: n_4544 <=  n_4545  AND n_4546;
delay_3861: n_4545  <= TRANSPORT a_LC6_F20  ;
delay_3862: n_4546  <= TRANSPORT a_LC4_F10  ;
and2_3863: n_4547 <=  n_4548  AND n_4549;
delay_3864: n_4548  <= TRANSPORT a_N757  ;
delay_3865: n_4549  <= TRANSPORT a_LC6_F20  ;
and2_3866: n_4550 <=  n_4551  AND n_4552;
delay_3867: n_4551  <= TRANSPORT a_N757  ;
delay_3868: n_4552  <= TRANSPORT a_LC4_F10  ;
and1_3869: n_4553 <=  gnd;
delay_3870: a_LC4_F15  <= TRANSPORT a_EQ004  ;
xor2_3871: a_EQ004 <=  n_4556  XOR n_4563;
or2_3872: n_4556 <=  n_4557  OR n_4560;
and2_3873: n_4557 <=  n_4558  AND n_4559;
delay_3874: n_4558  <= TRANSPORT a_LC6_F15  ;
inv_3875: n_4559  <= TRANSPORT NOT a_LC5_D27  ;
and2_3876: n_4560 <=  n_4561  AND n_4562;
inv_3877: n_4561  <= TRANSPORT NOT a_LC6_F15  ;
delay_3878: n_4562  <= TRANSPORT a_LC5_D27  ;
and1_3879: n_4563 <=  gnd;
delay_3880: a_LC1_F15  <= TRANSPORT a_EQ015  ;
xor2_3881: a_EQ015 <=  n_4566  XOR n_4573;
or2_3882: n_4566 <=  n_4567  OR n_4570;
and2_3883: n_4567 <=  n_4568  AND n_4569;
delay_3884: n_4568  <= TRANSPORT a_N757  ;
delay_3885: n_4569  <= TRANSPORT a_LC4_F15  ;
and2_3886: n_4570 <=  n_4571  AND n_4572;
delay_3887: n_4571  <= TRANSPORT a_LC6_F15  ;
delay_3888: n_4572  <= TRANSPORT a_LC5_D27  ;
and1_3889: n_4573 <=  gnd;
delay_3890: a_LC2_F14  <= TRANSPORT a_EQ295  ;
xor2_3891: a_EQ295 <=  n_4576  XOR n_4598;
or4_3892: n_4576 <=  n_4577  OR n_4583  OR n_4588  OR n_4593;
and4_3893: n_4577 <=  n_4578  AND n_4579  AND n_4580  AND n_4581;
inv_3894: n_4578  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_3895: n_4579  <= TRANSPORT a_N2529  ;
inv_3896: n_4580  <= TRANSPORT NOT a_LC1_F15  ;
inv_3897: n_4581  <= TRANSPORT NOT a_SADDRESSOUT_F8_G  ;
and4_3898: n_4583 <=  n_4584  AND n_4585  AND n_4586  AND n_4587;
inv_3899: n_4584  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_3900: n_4585  <= TRANSPORT NOT a_N2529  ;
inv_3901: n_4586  <= TRANSPORT NOT a_LC1_F15  ;
delay_3902: n_4587  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and4_3903: n_4588 <=  n_4589  AND n_4590  AND n_4591  AND n_4592;
inv_3904: n_4589  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_3905: n_4590  <= TRANSPORT NOT a_N2529  ;
delay_3906: n_4591  <= TRANSPORT a_LC1_F15  ;
inv_3907: n_4592  <= TRANSPORT NOT a_SADDRESSOUT_F8_G  ;
and4_3908: n_4593 <=  n_4594  AND n_4595  AND n_4596  AND n_4597;
inv_3909: n_4594  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_3910: n_4595  <= TRANSPORT a_N2529  ;
delay_3911: n_4596  <= TRANSPORT a_LC1_F15  ;
delay_3912: n_4597  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and1_3913: n_4598 <=  gnd;
delay_3914: a_LC1_F14  <= TRANSPORT a_EQ713  ;
xor2_3915: a_EQ713 <=  n_4601  XOR n_4611;
or2_3916: n_4601 <=  n_4602  OR n_4606;
and3_3917: n_4602 <=  n_4603  AND n_4604  AND n_4605;
inv_3918: n_4603  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_3919: n_4604  <= TRANSPORT a_N2560_aNOT  ;
delay_3920: n_4605  <= TRANSPORT dbin(0)  ;
and3_3921: n_4606 <=  n_4607  AND n_4608  AND n_4609;
delay_3922: n_4607  <= TRANSPORT a_N2583_aNOT  ;
delay_3923: n_4608  <= TRANSPORT a_N2560_aNOT  ;
delay_3924: n_4609  <= TRANSPORT a_SCH2ADDRREG_F8_G  ;
and1_3925: n_4611 <=  gnd;
dff_3926: DFF_a8237

    PORT MAP ( D => a_EQ1003, CLK => a_SCH2ADDRREG_F8_G_aCLK, CLRN => a_SCH2ADDRREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F8_G);
inv_3927: a_SCH2ADDRREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3928: a_EQ1003 <=  n_4618  XOR n_4628;
or3_3929: n_4618 <=  n_4619  OR n_4622  OR n_4625;
and2_3930: n_4619 <=  n_4620  AND n_4621;
inv_3931: n_4620  <= TRANSPORT NOT a_N2527  ;
delay_3932: n_4621  <= TRANSPORT a_LC2_F14  ;
and2_3933: n_4622 <=  n_4623  AND n_4624;
inv_3934: n_4623  <= TRANSPORT NOT a_N2527  ;
delay_3935: n_4624  <= TRANSPORT a_LC1_F14  ;
and2_3936: n_4625 <=  n_4626  AND n_4627;
delay_3937: n_4626  <= TRANSPORT a_SCH2BAROUT_F8_G  ;
delay_3938: n_4627  <= TRANSPORT a_N2527  ;
and1_3939: n_4628 <=  gnd;
delay_3940: n_4629  <= TRANSPORT clk  ;
filter_3941: FILTER_a8237

    PORT MAP (IN1 => n_4629, Y => a_SCH2ADDRREG_F8_G_aCLK);
delay_3942: a_LC5_D1  <= TRANSPORT a_EQ223  ;
xor2_3943: a_EQ223 <=  n_4633  XOR n_4641;
or2_3944: n_4633 <=  n_4634  OR n_4637;
and2_3945: n_4634 <=  n_4635  AND n_4636;
inv_3946: n_4635  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_3947: n_4636  <= TRANSPORT dbin(0)  ;
and2_3948: n_4637 <=  n_4638  AND n_4639;
delay_3949: n_4638  <= TRANSPORT a_N2573_aNOT  ;
delay_3950: n_4639  <= TRANSPORT a_SCH3WRDCNTREG_F8_G  ;
and1_3951: n_4641 <=  gnd;
delay_3952: a_LC6_D17  <= TRANSPORT a_EQ027  ;
xor2_3953: a_EQ027 <=  n_4644  XOR n_4655;
or3_3954: n_4644 <=  n_4645  OR n_4648  OR n_4651;
and2_3955: n_4645 <=  n_4646  AND n_4647;
delay_3956: n_4646  <= TRANSPORT a_N3549  ;
inv_3957: n_4647  <= TRANSPORT NOT a_N3548  ;
and2_3958: n_4648 <=  n_4649  AND n_4650;
inv_3959: n_4649  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
inv_3960: n_4650  <= TRANSPORT NOT a_N3548  ;
and3_3961: n_4651 <=  n_4652  AND n_4653  AND n_4654;
delay_3962: n_4652  <= TRANSPORT a_LC8_F13_aNOT  ;
inv_3963: n_4653  <= TRANSPORT NOT a_N3549  ;
delay_3964: n_4654  <= TRANSPORT a_N3548  ;
and1_3965: n_4655 <=  gnd;
delay_3966: a_LC6_D1  <= TRANSPORT a_EQ224  ;
xor2_3967: a_EQ224 <=  n_4658  XOR n_4665;
or2_3968: n_4658 <=  n_4659  OR n_4662;
and2_3969: n_4659 <=  n_4660  AND n_4661;
delay_3970: n_4660  <= TRANSPORT a_N965  ;
delay_3971: n_4661  <= TRANSPORT a_LC5_D1  ;
and2_3972: n_4662 <=  n_4663  AND n_4664;
inv_3973: n_4663  <= TRANSPORT NOT a_N965  ;
inv_3974: n_4664  <= TRANSPORT NOT a_LC6_D17  ;
and1_3975: n_4665 <=  gnd;
dff_3976: DFF_a8237

    PORT MAP ( D => a_EQ1121, CLK => a_SCH3WRDCNTREG_F8_G_aCLK, CLRN => a_SCH3WRDCNTREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F8_G);
inv_3977: a_SCH3WRDCNTREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_3978: a_EQ1121 <=  n_4672  XOR n_4679;
or2_3979: n_4672 <=  n_4673  OR n_4676;
and2_3980: n_4673 <=  n_4674  AND n_4675;
delay_3981: n_4674  <= TRANSPORT a_SCH3BWORDOUT_F8_G  ;
delay_3982: n_4675  <= TRANSPORT a_N2528  ;
and2_3983: n_4676 <=  n_4677  AND n_4678;
inv_3984: n_4677  <= TRANSPORT NOT a_N2528  ;
delay_3985: n_4678  <= TRANSPORT a_LC6_D1  ;
and1_3986: n_4679 <=  gnd;
delay_3987: n_4680  <= TRANSPORT clk  ;
filter_3988: FILTER_a8237

    PORT MAP (IN1 => n_4680, Y => a_SCH3WRDCNTREG_F8_G_aCLK);
delay_3989: a_N2548  <= TRANSPORT a_EQ605  ;
xor2_3990: a_EQ605 <=  n_4684  XOR n_4706;
or5_3991: n_4684 <=  n_4685  OR n_4689  OR n_4693  OR n_4696  OR n_4701;
and3_3992: n_4685 <=  n_4686  AND n_4687  AND n_4688;
delay_3993: n_4686  <= TRANSPORT a_N2529  ;
delay_3994: n_4687  <= TRANSPORT a_LC1_F15  ;
delay_3995: n_4688  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and3_3996: n_4689 <=  n_4690  AND n_4691  AND n_4692;
inv_3997: n_4690  <= TRANSPORT NOT a_N2529  ;
inv_3998: n_4691  <= TRANSPORT NOT a_LC1_F15  ;
delay_3999: n_4692  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and2_4000: n_4693 <=  n_4694  AND n_4695;
inv_4001: n_4694  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_4002: n_4695  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and4_4003: n_4696 <=  n_4697  AND n_4698  AND n_4699  AND n_4700;
inv_4004: n_4697  <= TRANSPORT NOT a_N2529  ;
delay_4005: n_4698  <= TRANSPORT a_N2530_aNOT  ;
delay_4006: n_4699  <= TRANSPORT a_LC1_F15  ;
inv_4007: n_4700  <= TRANSPORT NOT a_SADDRESSOUT_F8_G  ;
and4_4008: n_4701 <=  n_4702  AND n_4703  AND n_4704  AND n_4705;
delay_4009: n_4702  <= TRANSPORT a_N2529  ;
delay_4010: n_4703  <= TRANSPORT a_N2530_aNOT  ;
inv_4011: n_4704  <= TRANSPORT NOT a_LC1_F15  ;
inv_4012: n_4705  <= TRANSPORT NOT a_SADDRESSOUT_F8_G  ;
and1_4013: n_4706 <=  gnd;
delay_4014: a_LC1_F7  <= TRANSPORT a_EQ659  ;
xor2_4015: a_EQ659 <=  n_4709  XOR n_4717;
or2_4016: n_4709 <=  n_4710  OR n_4713;
and2_4017: n_4710 <=  n_4711  AND n_4712;
inv_4018: n_4711  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_4019: n_4712  <= TRANSPORT dbin(0)  ;
and2_4020: n_4713 <=  n_4714  AND n_4715;
delay_4021: n_4714  <= TRANSPORT a_N2587_aNOT  ;
delay_4022: n_4715  <= TRANSPORT a_SCH0ADDRREG_F8_G  ;
and1_4023: n_4717 <=  gnd;
delay_4024: a_LC2_F7  <= TRANSPORT a_EQ660  ;
xor2_4025: a_EQ660 <=  n_4720  XOR n_4727;
or2_4026: n_4720 <=  n_4721  OR n_4724;
and2_4027: n_4721 <=  n_4722  AND n_4723;
inv_4028: n_4722  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_4029: n_4723  <= TRANSPORT a_N2548  ;
and2_4030: n_4724 <=  n_4725  AND n_4726;
delay_4031: n_4725  <= TRANSPORT a_N2558_aNOT  ;
delay_4032: n_4726  <= TRANSPORT a_LC1_F7  ;
and1_4033: n_4727 <=  gnd;
dff_4034: DFF_a8237

    PORT MAP ( D => a_EQ875, CLK => a_SCH0ADDRREG_F8_G_aCLK, CLRN => a_SCH0ADDRREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F8_G);
inv_4035: a_SCH0ADDRREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4036: a_EQ875 <=  n_4734  XOR n_4741;
or2_4037: n_4734 <=  n_4735  OR n_4738;
and2_4038: n_4735 <=  n_4736  AND n_4737;
inv_4039: n_4736  <= TRANSPORT NOT a_N2525  ;
delay_4040: n_4737  <= TRANSPORT a_LC2_F7  ;
and2_4041: n_4738 <=  n_4739  AND n_4740;
delay_4042: n_4739  <= TRANSPORT a_SCH0BAROUT_F8_G  ;
delay_4043: n_4740  <= TRANSPORT a_N2525  ;
and1_4044: n_4741 <=  gnd;
delay_4045: n_4742  <= TRANSPORT clk  ;
filter_4046: FILTER_a8237

    PORT MAP (IN1 => n_4742, Y => a_SCH0ADDRREG_F8_G_aCLK);
delay_4047: a_LC5_F12  <= TRANSPORT a_EQ330  ;
xor2_4048: a_EQ330 <=  n_4746  XOR n_4767;
or4_4049: n_4746 <=  n_4747  OR n_4752  OR n_4757  OR n_4762;
and4_4050: n_4747 <=  n_4748  AND n_4749  AND n_4750  AND n_4751;
inv_4051: n_4748  <= TRANSPORT NOT a_N965  ;
inv_4052: n_4749  <= TRANSPORT NOT a_N2529  ;
delay_4053: n_4750  <= TRANSPORT a_LC1_F15  ;
inv_4054: n_4751  <= TRANSPORT NOT a_SADDRESSOUT_F8_G  ;
and4_4055: n_4752 <=  n_4753  AND n_4754  AND n_4755  AND n_4756;
inv_4056: n_4753  <= TRANSPORT NOT a_N965  ;
delay_4057: n_4754  <= TRANSPORT a_N2529  ;
delay_4058: n_4755  <= TRANSPORT a_LC1_F15  ;
delay_4059: n_4756  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and4_4060: n_4757 <=  n_4758  AND n_4759  AND n_4760  AND n_4761;
inv_4061: n_4758  <= TRANSPORT NOT a_N965  ;
delay_4062: n_4759  <= TRANSPORT a_N2529  ;
inv_4063: n_4760  <= TRANSPORT NOT a_LC1_F15  ;
inv_4064: n_4761  <= TRANSPORT NOT a_SADDRESSOUT_F8_G  ;
and4_4065: n_4762 <=  n_4763  AND n_4764  AND n_4765  AND n_4766;
inv_4066: n_4763  <= TRANSPORT NOT a_N965  ;
inv_4067: n_4764  <= TRANSPORT NOT a_N2529  ;
inv_4068: n_4765  <= TRANSPORT NOT a_LC1_F15  ;
delay_4069: n_4766  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and1_4070: n_4767 <=  gnd;
delay_4071: a_LC2_F12  <= TRANSPORT a_EQ738  ;
xor2_4072: a_EQ738 <=  n_4770  XOR n_4780;
or2_4073: n_4770 <=  n_4771  OR n_4775;
and3_4074: n_4771 <=  n_4772  AND n_4773  AND n_4774;
inv_4075: n_4772  <= TRANSPORT NOT a_N2581_aNOT  ;
delay_4076: n_4773  <= TRANSPORT a_N965  ;
delay_4077: n_4774  <= TRANSPORT dbin(0)  ;
and3_4078: n_4775 <=  n_4776  AND n_4777  AND n_4778;
delay_4079: n_4776  <= TRANSPORT a_N2581_aNOT  ;
delay_4080: n_4777  <= TRANSPORT a_N965  ;
delay_4081: n_4778  <= TRANSPORT a_SCH3ADDRREG_F8_G  ;
and1_4082: n_4780 <=  gnd;
dff_4083: DFF_a8237

    PORT MAP ( D => a_EQ1067, CLK => a_SCH3ADDRREG_F8_G_aCLK, CLRN => a_SCH3ADDRREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F8_G);
inv_4084: a_SCH3ADDRREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4085: a_EQ1067 <=  n_4787  XOR n_4797;
or3_4086: n_4787 <=  n_4788  OR n_4791  OR n_4794;
and2_4087: n_4788 <=  n_4789  AND n_4790;
inv_4088: n_4789  <= TRANSPORT NOT a_N2528  ;
delay_4089: n_4790  <= TRANSPORT a_LC5_F12  ;
and2_4090: n_4791 <=  n_4792  AND n_4793;
inv_4091: n_4792  <= TRANSPORT NOT a_N2528  ;
delay_4092: n_4793  <= TRANSPORT a_LC2_F12  ;
and2_4093: n_4794 <=  n_4795  AND n_4796;
delay_4094: n_4795  <= TRANSPORT a_SCH3BAROUT_F8_G  ;
delay_4095: n_4796  <= TRANSPORT a_N2528  ;
and1_4096: n_4797 <=  gnd;
delay_4097: n_4798  <= TRANSPORT clk  ;
filter_4098: FILTER_a8237

    PORT MAP (IN1 => n_4798, Y => a_SCH3ADDRREG_F8_G_aCLK);
delay_4099: a_LC6_D10  <= TRANSPORT a_EQ432  ;
xor2_4100: a_EQ432 <=  n_4802  XOR n_4814;
or3_4101: n_4802 <=  n_4803  OR n_4807  OR n_4811;
and3_4102: n_4803 <=  n_4804  AND n_4805  AND n_4806;
inv_4103: n_4804  <= TRANSPORT NOT a_LC3_D22  ;
inv_4104: n_4805  <= TRANSPORT NOT a_N2353  ;
delay_4105: n_4806  <= TRANSPORT dbin(0)  ;
and2_4106: n_4807 <=  n_4808  AND n_4809;
delay_4107: n_4808  <= TRANSPORT a_N2353  ;
delay_4108: n_4809  <= TRANSPORT a_SCH0WRDCNTREG_F8_G  ;
and2_4109: n_4811 <=  n_4812  AND n_4813;
delay_4110: n_4812  <= TRANSPORT a_LC3_D22  ;
delay_4111: n_4813  <= TRANSPORT a_SCH0WRDCNTREG_F8_G  ;
and1_4112: n_4814 <=  gnd;
delay_4113: a_LC8_D10  <= TRANSPORT a_EQ433  ;
xor2_4114: a_EQ433 <=  n_4817  XOR n_4824;
or2_4115: n_4817 <=  n_4818  OR n_4821;
and2_4116: n_4818 <=  n_4819  AND n_4820;
inv_4117: n_4819  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_4118: n_4820  <= TRANSPORT NOT a_LC6_D17  ;
and2_4119: n_4821 <=  n_4822  AND n_4823;
delay_4120: n_4822  <= TRANSPORT a_N2558_aNOT  ;
delay_4121: n_4823  <= TRANSPORT a_LC6_D10  ;
and1_4122: n_4824 <=  gnd;
dff_4123: DFF_a8237

    PORT MAP ( D => a_EQ929, CLK => a_SCH0WRDCNTREG_F8_G_aCLK, CLRN => a_SCH0WRDCNTREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F8_G);
inv_4124: a_SCH0WRDCNTREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4125: a_EQ929 <=  n_4831  XOR n_4838;
or2_4126: n_4831 <=  n_4832  OR n_4835;
and2_4127: n_4832 <=  n_4833  AND n_4834;
inv_4128: n_4833  <= TRANSPORT NOT a_N2525  ;
delay_4129: n_4834  <= TRANSPORT a_LC8_D10  ;
and2_4130: n_4835 <=  n_4836  AND n_4837;
delay_4131: n_4836  <= TRANSPORT a_SCH0BWORDOUT_F8_G  ;
delay_4132: n_4837  <= TRANSPORT a_N2525  ;
and1_4133: n_4838 <=  gnd;
delay_4134: n_4839  <= TRANSPORT clk  ;
filter_4135: FILTER_a8237

    PORT MAP (IN1 => n_4839, Y => a_SCH0WRDCNTREG_F8_G_aCLK);
delay_4136: a_N1553  <= TRANSPORT a_N1553_aIN  ;
xor2_4137: a_N1553_aIN <=  n_4843  XOR n_4847;
or1_4138: n_4843 <=  n_4844;
and2_4139: n_4844 <=  n_4845  AND n_4846;
inv_4140: n_4845  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_4141: n_4846  <= TRANSPORT a_N2548  ;
and1_4142: n_4847 <=  gnd;
delay_4143: a_LC7_F18  <= TRANSPORT a_EQ460  ;
xor2_4144: a_EQ460 <=  n_4850  XOR n_4860;
or2_4145: n_4850 <=  n_4851  OR n_4855;
and3_4146: n_4851 <=  n_4852  AND n_4853  AND n_4854;
inv_4147: n_4852  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_4148: n_4853  <= TRANSPORT a_N2559_aNOT  ;
delay_4149: n_4854  <= TRANSPORT dbin(0)  ;
and3_4150: n_4855 <=  n_4856  AND n_4857  AND n_4858;
delay_4151: n_4856  <= TRANSPORT a_N2585_aNOT  ;
delay_4152: n_4857  <= TRANSPORT a_N2559_aNOT  ;
delay_4153: n_4858  <= TRANSPORT a_SCH1ADDRREG_F8_G  ;
and1_4154: n_4860 <=  gnd;
dff_4155: DFF_a8237

    PORT MAP ( D => a_EQ939, CLK => a_SCH1ADDRREG_F8_G_aCLK, CLRN => a_SCH1ADDRREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F8_G);
inv_4156: a_SCH1ADDRREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4157: a_EQ939 <=  n_4867  XOR n_4877;
or3_4158: n_4867 <=  n_4868  OR n_4871  OR n_4874;
and2_4159: n_4868 <=  n_4869  AND n_4870;
inv_4160: n_4869  <= TRANSPORT NOT a_N2526  ;
delay_4161: n_4870  <= TRANSPORT a_N1553  ;
and2_4162: n_4871 <=  n_4872  AND n_4873;
inv_4163: n_4872  <= TRANSPORT NOT a_N2526  ;
delay_4164: n_4873  <= TRANSPORT a_LC7_F18  ;
and2_4165: n_4874 <=  n_4875  AND n_4876;
delay_4166: n_4875  <= TRANSPORT a_SCH1BAROUT_F8_G  ;
delay_4167: n_4876  <= TRANSPORT a_N2526  ;
and1_4168: n_4877 <=  gnd;
delay_4169: n_4878  <= TRANSPORT clk  ;
filter_4170: FILTER_a8237

    PORT MAP (IN1 => n_4878, Y => a_SCH1ADDRREG_F8_G_aCLK);
delay_4171: a_N689_aNOT  <= TRANSPORT a_EQ284  ;
xor2_4172: a_EQ284 <=  n_4882  XOR n_4894;
or3_4173: n_4882 <=  n_4883  OR n_4887  OR n_4891;
and3_4174: n_4883 <=  n_4884  AND n_4885  AND n_4886;
inv_4175: n_4884  <= TRANSPORT NOT a_LC3_D22  ;
inv_4176: n_4885  <= TRANSPORT NOT a_N62_aNOT  ;
delay_4177: n_4886  <= TRANSPORT dbin(0)  ;
and2_4178: n_4887 <=  n_4888  AND n_4889;
delay_4179: n_4888  <= TRANSPORT a_N62_aNOT  ;
delay_4180: n_4889  <= TRANSPORT a_SCH2WRDCNTREG_F8_G  ;
and2_4181: n_4891 <=  n_4892  AND n_4893;
delay_4182: n_4892  <= TRANSPORT a_LC3_D22  ;
delay_4183: n_4893  <= TRANSPORT a_SCH2WRDCNTREG_F8_G  ;
and1_4184: n_4894 <=  gnd;
delay_4185: a_LC3_D7  <= TRANSPORT a_EQ805  ;
xor2_4186: a_EQ805 <=  n_4897  XOR n_4904;
or2_4187: n_4897 <=  n_4898  OR n_4901;
and2_4188: n_4898 <=  n_4899  AND n_4900;
delay_4189: n_4899  <= TRANSPORT a_N2560_aNOT  ;
delay_4190: n_4900  <= TRANSPORT a_N689_aNOT  ;
and2_4191: n_4901 <=  n_4902  AND n_4903;
inv_4192: n_4902  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_4193: n_4903  <= TRANSPORT NOT a_LC6_D17  ;
and1_4194: n_4904 <=  gnd;
dff_4195: DFF_a8237

    PORT MAP ( D => a_EQ1057, CLK => a_SCH2WRDCNTREG_F8_G_aCLK, CLRN => a_SCH2WRDCNTREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F8_G);
inv_4196: a_SCH2WRDCNTREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4197: a_EQ1057 <=  n_4911  XOR n_4918;
or2_4198: n_4911 <=  n_4912  OR n_4915;
and2_4199: n_4912 <=  n_4913  AND n_4914;
inv_4200: n_4913  <= TRANSPORT NOT a_N2527  ;
delay_4201: n_4914  <= TRANSPORT a_LC3_D7  ;
and2_4202: n_4915 <=  n_4916  AND n_4917;
delay_4203: n_4916  <= TRANSPORT a_SCH2BWORDOUT_F8_G  ;
delay_4204: n_4917  <= TRANSPORT a_N2527  ;
and1_4205: n_4918 <=  gnd;
delay_4206: n_4919  <= TRANSPORT clk  ;
filter_4207: FILTER_a8237

    PORT MAP (IN1 => n_4919, Y => a_SCH2WRDCNTREG_F8_G_aCLK);
delay_4208: a_N357_aNOT  <= TRANSPORT a_EQ236  ;
xor2_4209: a_EQ236 <=  n_4923  XOR n_4931;
or2_4210: n_4923 <=  n_4924  OR n_4927;
and2_4211: n_4924 <=  n_4925  AND n_4926;
inv_4212: n_4925  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_4213: n_4926  <= TRANSPORT dbin(0)  ;
and2_4214: n_4927 <=  n_4928  AND n_4929;
delay_4215: n_4928  <= TRANSPORT a_N2577_aNOT  ;
delay_4216: n_4929  <= TRANSPORT a_SCH1WRDCNTREG_F8_G  ;
and1_4217: n_4931 <=  gnd;
delay_4218: a_LC3_D1  <= TRANSPORT a_EQ783  ;
xor2_4219: a_EQ783 <=  n_4934  XOR n_4941;
or2_4220: n_4934 <=  n_4935  OR n_4938;
and2_4221: n_4935 <=  n_4936  AND n_4937;
inv_4222: n_4936  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_4223: n_4937  <= TRANSPORT NOT a_LC6_D17  ;
and2_4224: n_4938 <=  n_4939  AND n_4940;
delay_4225: n_4939  <= TRANSPORT a_N2559_aNOT  ;
delay_4226: n_4940  <= TRANSPORT a_N357_aNOT  ;
and1_4227: n_4941 <=  gnd;
dff_4228: DFF_a8237

    PORT MAP ( D => a_EQ993, CLK => a_SCH1WRDCNTREG_F8_G_aCLK, CLRN => a_SCH1WRDCNTREG_F8_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F8_G);
inv_4229: a_SCH1WRDCNTREG_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4230: a_EQ993 <=  n_4948  XOR n_4955;
or2_4231: n_4948 <=  n_4949  OR n_4952;
and2_4232: n_4949 <=  n_4950  AND n_4951;
inv_4233: n_4950  <= TRANSPORT NOT a_N2526  ;
delay_4234: n_4951  <= TRANSPORT a_LC3_D1  ;
and2_4235: n_4952 <=  n_4953  AND n_4954;
delay_4236: n_4953  <= TRANSPORT a_SCH1BWORDOUT_F8_G  ;
delay_4237: n_4954  <= TRANSPORT a_N2526  ;
and1_4238: n_4955 <=  gnd;
delay_4239: n_4956  <= TRANSPORT clk  ;
filter_4240: FILTER_a8237

    PORT MAP (IN1 => n_4956, Y => a_SCH1WRDCNTREG_F8_G_aCLK);
delay_4241: a_LC3_D2  <= TRANSPORT a_EQ833  ;
xor2_4242: a_EQ833 <=  n_4960  XOR n_4969;
or2_4243: n_4960 <=  n_4961  OR n_4965;
and3_4244: n_4961 <=  n_4962  AND n_4963  AND n_4964;
inv_4245: n_4962  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_4246: n_4963  <= TRANSPORT a_N1095  ;
delay_4247: n_4964  <= TRANSPORT dbin(0)  ;
and3_4248: n_4965 <=  n_4966  AND n_4967  AND n_4968;
delay_4249: n_4966  <= TRANSPORT a_N2572_aNOT  ;
delay_4250: n_4967  <= TRANSPORT a_N1095  ;
delay_4251: n_4968  <= TRANSPORT a_SCH3WRDCNTREG_F0_G  ;
and1_4252: n_4969 <=  gnd;
delay_4253: a_N1033_aNOT  <= TRANSPORT a_N1033_aNOT_aIN  ;
xor2_4254: a_N1033_aNOT_aIN <=  n_4972  XOR n_4976;
or1_4255: n_4972 <=  n_4973;
and2_4256: n_4973 <=  n_4974  AND n_4975;
inv_4257: n_4974  <= TRANSPORT NOT a_N3556  ;
delay_4258: n_4975  <= TRANSPORT a_N1094  ;
and1_4259: n_4976 <=  gnd;
dff_4260: DFF_a8237

    PORT MAP ( D => a_EQ1113, CLK => a_SCH3WRDCNTREG_F0_G_aCLK, CLRN => a_SCH3WRDCNTREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F0_G);
inv_4261: a_SCH3WRDCNTREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4262: a_EQ1113 <=  n_4983  XOR n_4991;
or3_4263: n_4983 <=  n_4984  OR n_4986  OR n_4988;
and1_4264: n_4984 <=  n_4985;
delay_4265: n_4985  <= TRANSPORT a_LC3_D2  ;
and1_4266: n_4986 <=  n_4987;
delay_4267: n_4987  <= TRANSPORT a_N1033_aNOT  ;
and2_4268: n_4988 <=  n_4989  AND n_4990;
delay_4269: n_4989  <= TRANSPORT a_SCH3BWORDOUT_F0_G  ;
delay_4270: n_4990  <= TRANSPORT a_N2528  ;
and1_4271: n_4991 <=  gnd;
delay_4272: n_4992  <= TRANSPORT clk  ;
filter_4273: FILTER_a8237

    PORT MAP (IN1 => n_4992, Y => a_SCH3WRDCNTREG_F0_G_aCLK);
delay_4274: a_N241_aNOT  <= TRANSPORT a_EQ220  ;
xor2_4275: a_EQ220 <=  n_4996  XOR n_5003;
or2_4276: n_4996 <=  n_4997  OR n_5000;
and2_4277: n_4997 <=  n_4998  AND n_4999;
inv_4278: n_4998  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_4279: n_4999  <= TRANSPORT dbin(0)  ;
and2_4280: n_5000 <=  n_5001  AND n_5002;
delay_4281: n_5001  <= TRANSPORT a_N2578_aNOT  ;
delay_4282: n_5002  <= TRANSPORT a_SCH0WRDCNTREG_F0_G  ;
and1_4283: n_5003 <=  gnd;
delay_4284: a_LC2_D16  <= TRANSPORT a_EQ773  ;
xor2_4285: a_EQ773 <=  n_5006  XOR n_5013;
or2_4286: n_5006 <=  n_5007  OR n_5010;
and2_4287: n_5007 <=  n_5008  AND n_5009;
inv_4288: n_5008  <= TRANSPORT NOT a_N3556  ;
inv_4289: n_5009  <= TRANSPORT NOT a_N2558_aNOT  ;
and2_4290: n_5010 <=  n_5011  AND n_5012;
delay_4291: n_5011  <= TRANSPORT a_N2558_aNOT  ;
delay_4292: n_5012  <= TRANSPORT a_N241_aNOT  ;
and1_4293: n_5013 <=  gnd;
dff_4294: DFF_a8237

    PORT MAP ( D => a_EQ921, CLK => a_SCH0WRDCNTREG_F0_G_aCLK, CLRN => a_SCH0WRDCNTREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F0_G);
inv_4295: a_SCH0WRDCNTREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4296: a_EQ921 <=  n_5020  XOR n_5027;
or2_4297: n_5020 <=  n_5021  OR n_5024;
and2_4298: n_5021 <=  n_5022  AND n_5023;
inv_4299: n_5022  <= TRANSPORT NOT a_N2525  ;
delay_4300: n_5023  <= TRANSPORT a_LC2_D16  ;
and2_4301: n_5024 <=  n_5025  AND n_5026;
delay_4302: n_5025  <= TRANSPORT a_SCH0BWORDOUT_F0_G  ;
delay_4303: n_5026  <= TRANSPORT a_N2525  ;
and1_4304: n_5027 <=  gnd;
delay_4305: n_5028  <= TRANSPORT clk  ;
filter_4306: FILTER_a8237

    PORT MAP (IN1 => n_5028, Y => a_SCH0WRDCNTREG_F0_G_aCLK);
delay_4307: a_LC4_D20  <= TRANSPORT a_EQ813  ;
xor2_4308: a_EQ813 <=  n_5032  XOR n_5041;
or2_4309: n_5032 <=  n_5033  OR n_5037;
and3_4310: n_5033 <=  n_5034  AND n_5035  AND n_5036;
inv_4311: n_5034  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_4312: n_5035  <= TRANSPORT a_N756  ;
delay_4313: n_5036  <= TRANSPORT dbin(0)  ;
and3_4314: n_5037 <=  n_5038  AND n_5039  AND n_5040;
delay_4315: n_5038  <= TRANSPORT a_N2574_aNOT  ;
delay_4316: n_5039  <= TRANSPORT a_N756  ;
delay_4317: n_5040  <= TRANSPORT a_SCH2WRDCNTREG_F0_G  ;
and1_4318: n_5041 <=  gnd;
delay_4319: a_N805  <= TRANSPORT a_N805_aIN  ;
xor2_4320: a_N805_aIN <=  n_5044  XOR n_5048;
or1_4321: n_5044 <=  n_5045;
and2_4322: n_5045 <=  n_5046  AND n_5047;
inv_4323: n_5046  <= TRANSPORT NOT a_N3556  ;
delay_4324: n_5047  <= TRANSPORT a_N858  ;
and1_4325: n_5048 <=  gnd;
dff_4326: DFF_a8237

    PORT MAP ( D => a_EQ1049, CLK => a_SCH2WRDCNTREG_F0_G_aCLK, CLRN => a_SCH2WRDCNTREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F0_G);
inv_4327: a_SCH2WRDCNTREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4328: a_EQ1049 <=  n_5055  XOR n_5063;
or3_4329: n_5055 <=  n_5056  OR n_5058  OR n_5060;
and1_4330: n_5056 <=  n_5057;
delay_4331: n_5057  <= TRANSPORT a_LC4_D20  ;
and1_4332: n_5058 <=  n_5059;
delay_4333: n_5059  <= TRANSPORT a_N805  ;
and2_4334: n_5060 <=  n_5061  AND n_5062;
delay_4335: n_5061  <= TRANSPORT a_SCH2BWORDOUT_F0_G  ;
delay_4336: n_5062  <= TRANSPORT a_N2527  ;
and1_4337: n_5063 <=  gnd;
delay_4338: n_5064  <= TRANSPORT clk  ;
filter_4339: FILTER_a8237

    PORT MAP (IN1 => n_5064, Y => a_SCH2WRDCNTREG_F0_G_aCLK);
delay_4340: a_LC7_D16  <= TRANSPORT a_EQ794  ;
xor2_4341: a_EQ794 <=  n_5068  XOR n_5076;
or2_4342: n_5068 <=  n_5069  OR n_5072;
and2_4343: n_5069 <=  n_5070  AND n_5071;
delay_4344: n_5070  <= TRANSPORT a_LC7_D26  ;
delay_4345: n_5071  <= TRANSPORT a_SCH1WRDCNTREG_F0_G  ;
and2_4346: n_5072 <=  n_5073  AND n_5075;
delay_4347: n_5073  <= TRANSPORT a_SCH1BWORDOUT_F0_G  ;
delay_4348: n_5075  <= TRANSPORT a_N2526  ;
and1_4349: n_5076 <=  gnd;
delay_4350: a_N435  <= TRANSPORT a_N435_aIN  ;
xor2_4351: a_N435_aIN <=  n_5079  XOR n_5084;
or1_4352: n_5079 <=  n_5080;
and3_4353: n_5080 <=  n_5081  AND n_5082  AND n_5083;
inv_4354: n_5081  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_4355: n_5082  <= TRANSPORT a_N2595  ;
delay_4356: n_5083  <= TRANSPORT dbin(0)  ;
and1_4357: n_5084 <=  gnd;
dff_4358: DFF_a8237

    PORT MAP ( D => a_EQ985, CLK => a_SCH1WRDCNTREG_F0_G_aCLK, CLRN => a_SCH1WRDCNTREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F0_G);
inv_4359: a_SCH1WRDCNTREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4360: a_EQ985 <=  n_5091  XOR n_5099;
or3_4361: n_5091 <=  n_5092  OR n_5094  OR n_5096;
and1_4362: n_5092 <=  n_5093;
delay_4363: n_5093  <= TRANSPORT a_LC7_D16  ;
and1_4364: n_5094 <=  n_5095;
delay_4365: n_5095  <= TRANSPORT a_N435  ;
and2_4366: n_5096 <=  n_5097  AND n_5098;
inv_4367: n_5097  <= TRANSPORT NOT a_N3556  ;
delay_4368: n_5098  <= TRANSPORT a_N460  ;
and1_4369: n_5099 <=  gnd;
delay_4370: n_5100  <= TRANSPORT clk  ;
filter_4371: FILTER_a8237

    PORT MAP (IN1 => n_5100, Y => a_SCH1WRDCNTREG_F0_G_aCLK);
delay_4372: a_LC1_F10  <= TRANSPORT a_EQ014  ;
xor2_4373: a_EQ014 <=  n_5104  XOR n_5114;
or3_4374: n_5104 <=  n_5105  OR n_5108  OR n_5111;
and2_4375: n_5105 <=  n_5106  AND n_5107;
delay_4376: n_5106  <= TRANSPORT a_LC1_F15  ;
delay_4377: n_5107  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and2_4378: n_5108 <=  n_5109  AND n_5110;
delay_4379: n_5109  <= TRANSPORT a_N757  ;
delay_4380: n_5110  <= TRANSPORT a_LC1_F15  ;
and2_4381: n_5111 <=  n_5112  AND n_5113;
delay_4382: n_5112  <= TRANSPORT a_N757  ;
delay_4383: n_5113  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and1_4384: n_5114 <=  gnd;
delay_4385: a_LC3_A2  <= TRANSPORT a_EQ005  ;
xor2_4386: a_EQ005 <=  n_5117  XOR n_5125;
or2_4387: n_5117 <=  n_5118  OR n_5122;
and2_4388: n_5118 <=  n_5119  AND n_5120;
delay_4389: n_5119  <= TRANSPORT a_LC1_F10  ;
inv_4390: n_5120  <= TRANSPORT NOT a_SADDRESSOUT_F9_G  ;
and2_4391: n_5122 <=  n_5123  AND n_5124;
inv_4392: n_5123  <= TRANSPORT NOT a_LC1_F10  ;
delay_4393: n_5124  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
and1_4394: n_5125 <=  gnd;
delay_4395: a_LC4_A15  <= TRANSPORT a_EQ736  ;
xor2_4396: a_EQ736 <=  n_5128  XOR n_5140;
or3_4397: n_5128 <=  n_5129  OR n_5133  OR n_5137;
and3_4398: n_5129 <=  n_5130  AND n_5131  AND n_5132;
inv_4399: n_5130  <= TRANSPORT NOT a_LC3_D22  ;
inv_4400: n_5131  <= TRANSPORT NOT a_N2348  ;
delay_4401: n_5132  <= TRANSPORT dbin(1)  ;
and2_4402: n_5133 <=  n_5134  AND n_5135;
delay_4403: n_5134  <= TRANSPORT a_N2348  ;
delay_4404: n_5135  <= TRANSPORT a_SCH3ADDRREG_F9_G  ;
and2_4405: n_5137 <=  n_5138  AND n_5139;
delay_4406: n_5138  <= TRANSPORT a_LC3_D22  ;
delay_4407: n_5139  <= TRANSPORT a_SCH3ADDRREG_F9_G  ;
and1_4408: n_5140 <=  gnd;
delay_4409: a_LC6_A15  <= TRANSPORT a_EQ737  ;
xor2_4410: a_EQ737 <=  n_5143  XOR n_5155;
or3_4411: n_5143 <=  n_5144  OR n_5148  OR n_5152;
and3_4412: n_5144 <=  n_5145  AND n_5146  AND n_5147;
inv_4413: n_5145  <= TRANSPORT NOT a_N965  ;
inv_4414: n_5146  <= TRANSPORT NOT a_N2529  ;
delay_4415: n_5147  <= TRANSPORT a_LC3_A2  ;
and3_4416: n_5148 <=  n_5149  AND n_5150  AND n_5151;
inv_4417: n_5149  <= TRANSPORT NOT a_N965  ;
delay_4418: n_5150  <= TRANSPORT a_N2529  ;
inv_4419: n_5151  <= TRANSPORT NOT a_LC3_A2  ;
and2_4420: n_5152 <=  n_5153  AND n_5154;
delay_4421: n_5153  <= TRANSPORT a_N965  ;
delay_4422: n_5154  <= TRANSPORT a_LC4_A15  ;
and1_4423: n_5155 <=  gnd;
dff_4424: DFF_a8237

    PORT MAP ( D => a_EQ1068, CLK => a_SCH3ADDRREG_F9_G_aCLK, CLRN => a_SCH3ADDRREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F9_G);
inv_4425: a_SCH3ADDRREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4426: a_EQ1068 <=  n_5162  XOR n_5169;
or2_4427: n_5162 <=  n_5163  OR n_5166;
and2_4428: n_5163 <=  n_5164  AND n_5165;
inv_4429: n_5164  <= TRANSPORT NOT a_N2528  ;
delay_4430: n_5165  <= TRANSPORT a_LC6_A15  ;
and2_4431: n_5166 <=  n_5167  AND n_5168;
delay_4432: n_5167  <= TRANSPORT a_SCH3BAROUT_F9_G  ;
delay_4433: n_5168  <= TRANSPORT a_N2528  ;
and1_4434: n_5169 <=  gnd;
delay_4435: n_5170  <= TRANSPORT clk  ;
filter_4436: FILTER_a8237

    PORT MAP (IN1 => n_5170, Y => a_SCH3ADDRREG_F9_G_aCLK);
delay_4437: a_LC4_A16  <= TRANSPORT a_EQ711  ;
xor2_4438: a_EQ711 <=  n_5174  XOR n_5182;
or2_4439: n_5174 <=  n_5175  OR n_5178;
and2_4440: n_5175 <=  n_5176  AND n_5177;
inv_4441: n_5176  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_4442: n_5177  <= TRANSPORT dbin(1)  ;
and2_4443: n_5178 <=  n_5179  AND n_5180;
delay_4444: n_5179  <= TRANSPORT a_N2583_aNOT  ;
delay_4445: n_5180  <= TRANSPORT a_SCH2ADDRREG_F9_G  ;
and1_4446: n_5182 <=  gnd;
delay_4447: a_LC6_A16  <= TRANSPORT a_EQ712  ;
xor2_4448: a_EQ712 <=  n_5185  XOR n_5197;
or3_4449: n_5185 <=  n_5186  OR n_5190  OR n_5194;
and3_4450: n_5186 <=  n_5187  AND n_5188  AND n_5189;
inv_4451: n_5187  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_4452: n_5188  <= TRANSPORT NOT a_N2529  ;
delay_4453: n_5189  <= TRANSPORT a_LC3_A2  ;
and3_4454: n_5190 <=  n_5191  AND n_5192  AND n_5193;
inv_4455: n_5191  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_4456: n_5192  <= TRANSPORT a_N2529  ;
inv_4457: n_5193  <= TRANSPORT NOT a_LC3_A2  ;
and2_4458: n_5194 <=  n_5195  AND n_5196;
delay_4459: n_5195  <= TRANSPORT a_N2560_aNOT  ;
delay_4460: n_5196  <= TRANSPORT a_LC4_A16  ;
and1_4461: n_5197 <=  gnd;
dff_4462: DFF_a8237

    PORT MAP ( D => a_EQ1004, CLK => a_SCH2ADDRREG_F9_G_aCLK, CLRN => a_SCH2ADDRREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F9_G);
inv_4463: a_SCH2ADDRREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4464: a_EQ1004 <=  n_5204  XOR n_5211;
or2_4465: n_5204 <=  n_5205  OR n_5208;
and2_4466: n_5205 <=  n_5206  AND n_5207;
inv_4467: n_5206  <= TRANSPORT NOT a_N2527  ;
delay_4468: n_5207  <= TRANSPORT a_LC6_A16  ;
and2_4469: n_5208 <=  n_5209  AND n_5210;
delay_4470: n_5209  <= TRANSPORT a_SCH2BAROUT_F9_G  ;
delay_4471: n_5210  <= TRANSPORT a_N2527  ;
and1_4472: n_5211 <=  gnd;
delay_4473: n_5212  <= TRANSPORT clk  ;
filter_4474: FILTER_a8237

    PORT MAP (IN1 => n_5212, Y => a_SCH2ADDRREG_F9_G_aCLK);
delay_4475: a_N2549  <= TRANSPORT a_EQ606  ;
xor2_4476: a_EQ606 <=  n_5216  XOR n_5228;
or3_4477: n_5216 <=  n_5217  OR n_5221  OR n_5225;
and3_4478: n_5217 <=  n_5218  AND n_5219  AND n_5220;
inv_4479: n_5218  <= TRANSPORT NOT a_N2529  ;
delay_4480: n_5219  <= TRANSPORT a_N2530_aNOT  ;
delay_4481: n_5220  <= TRANSPORT a_LC3_A2  ;
and3_4482: n_5221 <=  n_5222  AND n_5223  AND n_5224;
delay_4483: n_5222  <= TRANSPORT a_N2529  ;
delay_4484: n_5223  <= TRANSPORT a_N2530_aNOT  ;
inv_4485: n_5224  <= TRANSPORT NOT a_LC3_A2  ;
and2_4486: n_5225 <=  n_5226  AND n_5227;
inv_4487: n_5226  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_4488: n_5227  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
and1_4489: n_5228 <=  gnd;
delay_4490: a_LC4_A8  <= TRANSPORT a_EQ657  ;
xor2_4491: a_EQ657 <=  n_5231  XOR n_5243;
or3_4492: n_5231 <=  n_5232  OR n_5236  OR n_5240;
and3_4493: n_5232 <=  n_5233  AND n_5234  AND n_5235;
inv_4494: n_5233  <= TRANSPORT NOT a_LC3_D22  ;
delay_4495: n_5234  <= TRANSPORT a_N2354_aNOT  ;
delay_4496: n_5235  <= TRANSPORT dbin(1)  ;
and2_4497: n_5236 <=  n_5237  AND n_5238;
inv_4498: n_5237  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_4499: n_5238  <= TRANSPORT a_SCH0ADDRREG_F9_G  ;
and2_4500: n_5240 <=  n_5241  AND n_5242;
delay_4501: n_5241  <= TRANSPORT a_LC3_D22  ;
delay_4502: n_5242  <= TRANSPORT a_SCH0ADDRREG_F9_G  ;
and1_4503: n_5243 <=  gnd;
delay_4504: a_LC3_A8  <= TRANSPORT a_EQ658  ;
xor2_4505: a_EQ658 <=  n_5246  XOR n_5253;
or2_4506: n_5246 <=  n_5247  OR n_5250;
and2_4507: n_5247 <=  n_5248  AND n_5249;
inv_4508: n_5248  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_4509: n_5249  <= TRANSPORT a_N2549  ;
and2_4510: n_5250 <=  n_5251  AND n_5252;
delay_4511: n_5251  <= TRANSPORT a_N2558_aNOT  ;
delay_4512: n_5252  <= TRANSPORT a_LC4_A8  ;
and1_4513: n_5253 <=  gnd;
dff_4514: DFF_a8237

    PORT MAP ( D => a_EQ876, CLK => a_SCH0ADDRREG_F9_G_aCLK, CLRN => a_SCH0ADDRREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F9_G);
inv_4515: a_SCH0ADDRREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4516: a_EQ876 <=  n_5260  XOR n_5267;
or2_4517: n_5260 <=  n_5261  OR n_5264;
and2_4518: n_5261 <=  n_5262  AND n_5263;
inv_4519: n_5262  <= TRANSPORT NOT a_N2525  ;
delay_4520: n_5263  <= TRANSPORT a_LC3_A8  ;
and2_4521: n_5264 <=  n_5265  AND n_5266;
delay_4522: n_5265  <= TRANSPORT a_SCH0BAROUT_F9_G  ;
delay_4523: n_5266  <= TRANSPORT a_N2525  ;
and1_4524: n_5267 <=  gnd;
delay_4525: n_5268  <= TRANSPORT clk  ;
filter_4526: FILTER_a8237

    PORT MAP (IN1 => n_5268, Y => a_SCH0ADDRREG_F9_G_aCLK);
delay_4527: a_LC2_A12  <= TRANSPORT a_EQ683  ;
xor2_4528: a_EQ683 <=  n_5272  XOR n_5284;
or3_4529: n_5272 <=  n_5273  OR n_5277  OR n_5281;
and3_4530: n_5273 <=  n_5274  AND n_5275  AND n_5276;
inv_4531: n_5274  <= TRANSPORT NOT a_LC3_D22  ;
inv_4532: n_5275  <= TRANSPORT NOT a_N2352  ;
delay_4533: n_5276  <= TRANSPORT dbin(1)  ;
and2_4534: n_5277 <=  n_5278  AND n_5279;
delay_4535: n_5278  <= TRANSPORT a_N2352  ;
delay_4536: n_5279  <= TRANSPORT a_SCH1ADDRREG_F9_G  ;
and2_4537: n_5281 <=  n_5282  AND n_5283;
delay_4538: n_5282  <= TRANSPORT a_LC3_D22  ;
delay_4539: n_5283  <= TRANSPORT a_SCH1ADDRREG_F9_G  ;
and1_4540: n_5284 <=  gnd;
delay_4541: a_LC3_A12  <= TRANSPORT a_EQ684  ;
xor2_4542: a_EQ684 <=  n_5287  XOR n_5294;
or2_4543: n_5287 <=  n_5288  OR n_5291;
and2_4544: n_5288 <=  n_5289  AND n_5290;
inv_4545: n_5289  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_4546: n_5290  <= TRANSPORT a_N2549  ;
and2_4547: n_5291 <=  n_5292  AND n_5293;
delay_4548: n_5292  <= TRANSPORT a_N2559_aNOT  ;
delay_4549: n_5293  <= TRANSPORT a_LC2_A12  ;
and1_4550: n_5294 <=  gnd;
dff_4551: DFF_a8237

    PORT MAP ( D => a_EQ940, CLK => a_SCH1ADDRREG_F9_G_aCLK, CLRN => a_SCH1ADDRREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F9_G);
inv_4552: a_SCH1ADDRREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4553: a_EQ940 <=  n_5301  XOR n_5308;
or2_4554: n_5301 <=  n_5302  OR n_5305;
and2_4555: n_5302 <=  n_5303  AND n_5304;
inv_4556: n_5303  <= TRANSPORT NOT a_N2526  ;
delay_4557: n_5304  <= TRANSPORT a_LC3_A12  ;
and2_4558: n_5305 <=  n_5306  AND n_5307;
delay_4559: n_5306  <= TRANSPORT a_N2526  ;
delay_4560: n_5307  <= TRANSPORT a_SCH1BAROUT_F9_G  ;
and1_4561: n_5308 <=  gnd;
delay_4562: n_5309  <= TRANSPORT clk  ;
filter_4563: FILTER_a8237

    PORT MAP (IN1 => n_5309, Y => a_SCH1ADDRREG_F9_G_aCLK);
delay_4564: a_LC2_A21  <= TRANSPORT a_EQ824  ;
xor2_4565: a_EQ824 <=  n_5313  XOR n_5321;
or2_4566: n_5313 <=  n_5314  OR n_5317;
and2_4567: n_5314 <=  n_5315  AND n_5316;
inv_4568: n_5315  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_4569: n_5316  <= TRANSPORT dbin(1)  ;
and2_4570: n_5317 <=  n_5318  AND n_5319;
delay_4571: n_5318  <= TRANSPORT a_N2573_aNOT  ;
delay_4572: n_5319  <= TRANSPORT a_SCH3WRDCNTREG_F9_G  ;
and1_4573: n_5321 <=  gnd;
delay_4574: a_LC1_A21  <= TRANSPORT a_EQ825  ;
xor2_4575: a_EQ825 <=  n_5324  XOR n_5335;
or3_4576: n_5324 <=  n_5325  OR n_5329  OR n_5332;
and3_4577: n_5325 <=  n_5326  AND n_5327  AND n_5328;
delay_4578: n_5326  <= TRANSPORT a_N2557  ;
inv_4579: n_5327  <= TRANSPORT NOT a_N2377  ;
inv_4580: n_5328  <= TRANSPORT NOT a_LC1_A13  ;
and2_4581: n_5329 <=  n_5330  AND n_5331;
inv_4582: n_5330  <= TRANSPORT NOT a_N2557  ;
delay_4583: n_5331  <= TRANSPORT a_LC2_A21  ;
and2_4584: n_5332 <=  n_5333  AND n_5334;
delay_4585: n_5333  <= TRANSPORT a_N2377  ;
delay_4586: n_5334  <= TRANSPORT a_LC2_A21  ;
and1_4587: n_5335 <=  gnd;
dff_4588: DFF_a8237

    PORT MAP ( D => a_EQ1122, CLK => a_SCH3WRDCNTREG_F9_G_aCLK, CLRN => a_SCH3WRDCNTREG_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F9_G);
inv_4589: a_SCH3WRDCNTREG_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4590: a_EQ1122 <=  n_5342  XOR n_5349;
or2_4591: n_5342 <=  n_5343  OR n_5346;
and2_4592: n_5343 <=  n_5344  AND n_5345;
inv_4593: n_5344  <= TRANSPORT NOT a_N2528  ;
delay_4594: n_5345  <= TRANSPORT a_LC1_A21  ;
and2_4595: n_5346 <=  n_5347  AND n_5348;
delay_4596: n_5347  <= TRANSPORT a_N2528  ;
delay_4597: n_5348  <= TRANSPORT a_SCH3BWORDOUT_F9_G  ;
and1_4598: n_5349 <=  gnd;
delay_4599: n_5350  <= TRANSPORT clk  ;
filter_4600: FILTER_a8237

    PORT MAP (IN1 => n_5350, Y => a_SCH3WRDCNTREG_F9_G_aCLK);
delay_4601: a_N2367  <= TRANSPORT a_EQ563  ;
xor2_4602: a_EQ563 <=  n_5354  XOR n_5363;
or4_4603: n_5354 <=  n_5355  OR n_5357  OR n_5359  OR n_5361;
and1_4604: n_5355 <=  n_5356;
delay_4605: n_5356  <= TRANSPORT ain(2)  ;
and1_4606: n_5357 <=  n_5358;
delay_4607: n_5358  <= TRANSPORT ain(1)  ;
and1_4608: n_5359 <=  n_5360;
delay_4609: n_5360  <= TRANSPORT ain(0)  ;
and1_4610: n_5361 <=  n_5362;
inv_4611: n_5362  <= TRANSPORT NOT ain(3)  ;
and1_4612: n_5363 <=  gnd;
dff_4613: DFF_a8237

    PORT MAP ( D => a_N824_aD, CLK => a_N824_aCLK, CLRN => a_N824_aCLRN, PRN => vcc,
          Q => a_N824);
inv_4614: a_N824_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4615: a_N824_aD <=  n_5371  XOR n_5375;
or1_4616: n_5371 <=  n_5372;
and1_4617: n_5372 <=  n_5373;
delay_4618: n_5373  <= TRANSPORT niorin  ;
and1_4619: n_5375 <=  gnd;
delay_4620: n_5376  <= TRANSPORT clk  ;
filter_4621: FILTER_a8237

    PORT MAP (IN1 => n_5376, Y => a_N824_aCLK);
delay_4622: a_LC2_B15  <= TRANSPORT a_LC2_B15_aIN  ;
xor2_4623: a_LC2_B15_aIN <=  n_5380  XOR n_5386;
or1_4624: n_5380 <=  n_5381;
and3_4625: n_5381 <=  n_5382  AND n_5383  AND n_5384;
inv_4626: n_5382  <= TRANSPORT NOT a_N824  ;
delay_4627: n_5383  <= TRANSPORT niorin  ;
inv_4628: n_5384  <= TRANSPORT NOT ncs  ;
and1_4629: n_5386 <=  gnd;
delay_4630: a_N2592  <= TRANSPORT a_EQ643  ;
xor2_4631: a_EQ643 <=  n_5389  XOR n_5398;
or2_4632: n_5389 <=  n_5390  OR n_5394;
and3_4633: n_5390 <=  n_5391  AND n_5392  AND n_5393;
delay_4634: n_5391  <= TRANSPORT a_N2563_aNOT  ;
delay_4635: n_5392  <= TRANSPORT a_N2367  ;
inv_4636: n_5393  <= TRANSPORT NOT reset  ;
and3_4637: n_5394 <=  n_5395  AND n_5396  AND n_5397;
delay_4638: n_5395  <= TRANSPORT a_N2563_aNOT  ;
inv_4639: n_5396  <= TRANSPORT NOT a_LC2_B15  ;
inv_4640: n_5397  <= TRANSPORT NOT reset  ;
and1_4641: n_5398 <=  gnd;
delay_4642: a_N1523  <= TRANSPORT a_EQ457  ;
xor2_4643: a_EQ457 <=  n_5401  XOR n_5406;
or2_4644: n_5401 <=  n_5402  OR n_5404;
and1_4645: n_5402 <=  n_5403;
delay_4646: n_5403  <= TRANSPORT a_N2591  ;
and1_4647: n_5404 <=  n_5405;
inv_4648: n_5405  <= TRANSPORT NOT a_N88_aNOT  ;
and1_4649: n_5406 <=  gnd;
dff_4650: DFF_a8237

    PORT MAP ( D => a_EQ1178, CLK => a_STCSTATUS_F1_G_aCLK, CLRN => a_STCSTATUS_F1_G_aCLRN,
          PRN => vcc, Q => a_STCSTATUS_F1_G);
inv_4651: a_STCSTATUS_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4652: a_EQ1178 <=  n_5414  XOR n_5422;
or2_4653: n_5414 <=  n_5415  OR n_5418;
and2_4654: n_5415 <=  n_5416  AND n_5417;
delay_4655: n_5416  <= TRANSPORT a_N2592  ;
delay_4656: n_5417  <= TRANSPORT a_STCSTATUS_F1_G  ;
and3_4657: n_5418 <=  n_5419  AND n_5420  AND n_5421;
delay_4658: n_5419  <= TRANSPORT a_N57_aNOT  ;
delay_4659: n_5420  <= TRANSPORT a_N2592  ;
delay_4660: n_5421  <= TRANSPORT a_N1523  ;
and1_4661: n_5422 <=  gnd;
delay_4662: n_5423  <= TRANSPORT clk  ;
filter_4663: FILTER_a8237

    PORT MAP (IN1 => n_5423, Y => a_STCSTATUS_F1_G_aCLK);
delay_4664: a_LC5_C4  <= TRANSPORT a_EQ831  ;
xor2_4665: a_EQ831 <=  n_5427  XOR n_5436;
or2_4666: n_5427 <=  n_5428  OR n_5432;
and3_4667: n_5428 <=  n_5429  AND n_5430  AND n_5431;
inv_4668: n_5429  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_4669: n_5430  <= TRANSPORT a_N1095  ;
delay_4670: n_5431  <= TRANSPORT dbin(2)  ;
and3_4671: n_5432 <=  n_5433  AND n_5434  AND n_5435;
delay_4672: n_5433  <= TRANSPORT a_N2572_aNOT  ;
delay_4673: n_5434  <= TRANSPORT a_N1095  ;
delay_4674: n_5435  <= TRANSPORT a_SCH3WRDCNTREG_F2_G  ;
and1_4675: n_5436 <=  gnd;
delay_4676: a_N1047_aNOT  <= TRANSPORT a_N1047_aNOT_aIN  ;
xor2_4677: a_N1047_aNOT_aIN <=  n_5439  XOR n_5443;
or1_4678: n_5439 <=  n_5440;
and2_4679: n_5440 <=  n_5441  AND n_5442;
delay_4680: n_5441  <= TRANSPORT a_SCH3BWORDOUT_F2_G  ;
delay_4681: n_5442  <= TRANSPORT a_N2528  ;
and1_4682: n_5443 <=  gnd;
dff_4683: DFF_a8237

    PORT MAP ( D => a_EQ1115, CLK => a_SCH3WRDCNTREG_F2_G_aCLK, CLRN => a_SCH3WRDCNTREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F2_G);
inv_4684: a_SCH3WRDCNTREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4685: a_EQ1115 <=  n_5450  XOR n_5458;
or3_4686: n_5450 <=  n_5451  OR n_5453  OR n_5455;
and1_4687: n_5451 <=  n_5452;
delay_4688: n_5452  <= TRANSPORT a_LC5_C4  ;
and1_4689: n_5453 <=  n_5454;
delay_4690: n_5454  <= TRANSPORT a_N1047_aNOT  ;
and2_4691: n_5455 <=  n_5456  AND n_5457;
inv_4692: n_5456  <= TRANSPORT NOT a_LC1_C22  ;
delay_4693: n_5457  <= TRANSPORT a_N1094  ;
and1_4694: n_5458 <=  gnd;
delay_4695: n_5459  <= TRANSPORT clk  ;
filter_4696: FILTER_a8237

    PORT MAP (IN1 => n_5459, Y => a_SCH3WRDCNTREG_F2_G_aCLK);
delay_4697: a_LC1_D20  <= TRANSPORT a_EQ811  ;
xor2_4698: a_EQ811 <=  n_5463  XOR n_5472;
or2_4699: n_5463 <=  n_5464  OR n_5468;
and3_4700: n_5464 <=  n_5465  AND n_5466  AND n_5467;
inv_4701: n_5465  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_4702: n_5466  <= TRANSPORT a_N756  ;
delay_4703: n_5467  <= TRANSPORT dbin(2)  ;
and3_4704: n_5468 <=  n_5469  AND n_5470  AND n_5471;
delay_4705: n_5469  <= TRANSPORT a_N2574_aNOT  ;
delay_4706: n_5470  <= TRANSPORT a_N756  ;
delay_4707: n_5471  <= TRANSPORT a_SCH2WRDCNTREG_F2_G  ;
and1_4708: n_5472 <=  gnd;
delay_4709: a_N799  <= TRANSPORT a_N799_aIN  ;
xor2_4710: a_N799_aIN <=  n_5475  XOR n_5479;
or1_4711: n_5475 <=  n_5476;
and2_4712: n_5476 <=  n_5477  AND n_5478;
delay_4713: n_5477  <= TRANSPORT a_SCH2BWORDOUT_F2_G  ;
delay_4714: n_5478  <= TRANSPORT a_N2527  ;
and1_4715: n_5479 <=  gnd;
dff_4716: DFF_a8237

    PORT MAP ( D => a_EQ1051, CLK => a_SCH2WRDCNTREG_F2_G_aCLK, CLRN => a_SCH2WRDCNTREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F2_G);
inv_4717: a_SCH2WRDCNTREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4718: a_EQ1051 <=  n_5486  XOR n_5494;
or3_4719: n_5486 <=  n_5487  OR n_5489  OR n_5491;
and1_4720: n_5487 <=  n_5488;
delay_4721: n_5488  <= TRANSPORT a_LC1_D20  ;
and1_4722: n_5489 <=  n_5490;
delay_4723: n_5490  <= TRANSPORT a_N799  ;
and2_4724: n_5491 <=  n_5492  AND n_5493;
inv_4725: n_5492  <= TRANSPORT NOT a_LC1_C22  ;
delay_4726: n_5493  <= TRANSPORT a_N858  ;
and1_4727: n_5494 <=  gnd;
delay_4728: n_5495  <= TRANSPORT clk  ;
filter_4729: FILTER_a8237

    PORT MAP (IN1 => n_5495, Y => a_SCH2WRDCNTREG_F2_G_aCLK);
delay_4730: a_LC3_C3  <= TRANSPORT a_EQ769  ;
xor2_4731: a_EQ769 <=  n_5499  XOR n_5506;
or2_4732: n_5499 <=  n_5500  OR n_5503;
and2_4733: n_5500 <=  n_5501  AND n_5502;
inv_4734: n_5501  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_4735: n_5502  <= TRANSPORT dbin(2)  ;
and2_4736: n_5503 <=  n_5504  AND n_5505;
delay_4737: n_5504  <= TRANSPORT a_N2578_aNOT  ;
delay_4738: n_5505  <= TRANSPORT a_SCH0WRDCNTREG_F2_G  ;
and1_4739: n_5506 <=  gnd;
delay_4740: a_LC5_C3  <= TRANSPORT a_EQ770  ;
xor2_4741: a_EQ770 <=  n_5509  XOR n_5516;
or2_4742: n_5509 <=  n_5510  OR n_5513;
and2_4743: n_5510 <=  n_5511  AND n_5512;
inv_4744: n_5511  <= TRANSPORT NOT a_LC1_C22  ;
inv_4745: n_5512  <= TRANSPORT NOT a_N2558_aNOT  ;
and2_4746: n_5513 <=  n_5514  AND n_5515;
delay_4747: n_5514  <= TRANSPORT a_N2558_aNOT  ;
delay_4748: n_5515  <= TRANSPORT a_LC3_C3  ;
and1_4749: n_5516 <=  gnd;
dff_4750: DFF_a8237

    PORT MAP ( D => a_EQ923, CLK => a_SCH0WRDCNTREG_F2_G_aCLK, CLRN => a_SCH0WRDCNTREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F2_G);
inv_4751: a_SCH0WRDCNTREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4752: a_EQ923 <=  n_5523  XOR n_5530;
or2_4753: n_5523 <=  n_5524  OR n_5527;
and2_4754: n_5524 <=  n_5525  AND n_5526;
inv_4755: n_5525  <= TRANSPORT NOT a_N2525  ;
delay_4756: n_5526  <= TRANSPORT a_LC5_C3  ;
and2_4757: n_5527 <=  n_5528  AND n_5529;
delay_4758: n_5528  <= TRANSPORT a_N2525  ;
delay_4759: n_5529  <= TRANSPORT a_SCH0BWORDOUT_F2_G  ;
and1_4760: n_5530 <=  gnd;
delay_4761: n_5531  <= TRANSPORT clk  ;
filter_4762: FILTER_a8237

    PORT MAP (IN1 => n_5531, Y => a_SCH0WRDCNTREG_F2_G_aCLK);
delay_4763: a_LC3_D26  <= TRANSPORT a_EQ792  ;
xor2_4764: a_EQ792 <=  n_5535  XOR n_5543;
or2_4765: n_5535 <=  n_5536  OR n_5539;
and2_4766: n_5536 <=  n_5537  AND n_5538;
delay_4767: n_5537  <= TRANSPORT a_LC7_D26  ;
delay_4768: n_5538  <= TRANSPORT a_SCH1WRDCNTREG_F2_G  ;
and2_4769: n_5539 <=  n_5540  AND n_5542;
delay_4770: n_5540  <= TRANSPORT a_SCH1BWORDOUT_F2_G  ;
delay_4771: n_5542  <= TRANSPORT a_N2526  ;
and1_4772: n_5543 <=  gnd;
delay_4773: a_N434  <= TRANSPORT a_N434_aIN  ;
xor2_4774: a_N434_aIN <=  n_5546  XOR n_5552;
or1_4775: n_5546 <=  n_5547;
and4_4776: n_5547 <=  n_5548  AND n_5549  AND n_5550  AND n_5551;
inv_4777: n_5548  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_4778: n_5549  <= TRANSPORT a_N2559_aNOT  ;
inv_4779: n_5550  <= TRANSPORT NOT a_N2526  ;
delay_4780: n_5551  <= TRANSPORT dbin(2)  ;
and1_4781: n_5552 <=  gnd;
dff_4782: DFF_a8237

    PORT MAP ( D => a_EQ987, CLK => a_SCH1WRDCNTREG_F2_G_aCLK, CLRN => a_SCH1WRDCNTREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F2_G);
inv_4783: a_SCH1WRDCNTREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4784: a_EQ987 <=  n_5559  XOR n_5567;
or3_4785: n_5559 <=  n_5560  OR n_5562  OR n_5564;
and1_4786: n_5560 <=  n_5561;
delay_4787: n_5561  <= TRANSPORT a_LC3_D26  ;
and1_4788: n_5562 <=  n_5563;
delay_4789: n_5563  <= TRANSPORT a_N434  ;
and2_4790: n_5564 <=  n_5565  AND n_5566;
inv_4791: n_5565  <= TRANSPORT NOT a_LC1_C22  ;
delay_4792: n_5566  <= TRANSPORT a_N460  ;
and1_4793: n_5567 <=  gnd;
delay_4794: n_5568  <= TRANSPORT clk  ;
filter_4795: FILTER_a8237

    PORT MAP (IN1 => n_5568, Y => a_SCH1WRDCNTREG_F2_G_aCLK);
delay_4796: a_LC2_A9  <= TRANSPORT a_EQ006  ;
xor2_4797: a_EQ006 <=  n_5572  XOR n_5598;
or6_4798: n_5572 <=  n_5573  OR n_5578  OR n_5582  OR n_5586  OR n_5590  OR n_5594;
and3_4799: n_5573 <=  n_5574  AND n_5575  AND n_5576;
delay_4800: n_5574  <= TRANSPORT a_LC1_F10  ;
delay_4801: n_5575  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
inv_4802: n_5576  <= TRANSPORT NOT a_SADDRESSOUT_F10_G  ;
and3_4803: n_5578 <=  n_5579  AND n_5580  AND n_5581;
delay_4804: n_5579  <= TRANSPORT a_N757  ;
delay_4805: n_5580  <= TRANSPORT a_LC1_F10  ;
inv_4806: n_5581  <= TRANSPORT NOT a_SADDRESSOUT_F10_G  ;
and3_4807: n_5582 <=  n_5583  AND n_5584  AND n_5585;
delay_4808: n_5583  <= TRANSPORT a_N757  ;
delay_4809: n_5584  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
inv_4810: n_5585  <= TRANSPORT NOT a_SADDRESSOUT_F10_G  ;
and3_4811: n_5586 <=  n_5587  AND n_5588  AND n_5589;
inv_4812: n_5587  <= TRANSPORT NOT a_LC1_F10  ;
inv_4813: n_5588  <= TRANSPORT NOT a_SADDRESSOUT_F9_G  ;
delay_4814: n_5589  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and3_4815: n_5590 <=  n_5591  AND n_5592  AND n_5593;
inv_4816: n_5591  <= TRANSPORT NOT a_N757  ;
inv_4817: n_5592  <= TRANSPORT NOT a_SADDRESSOUT_F9_G  ;
delay_4818: n_5593  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and3_4819: n_5594 <=  n_5595  AND n_5596  AND n_5597;
inv_4820: n_5595  <= TRANSPORT NOT a_N757  ;
inv_4821: n_5596  <= TRANSPORT NOT a_LC1_F10  ;
delay_4822: n_5597  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and1_4823: n_5598 <=  gnd;
delay_4824: a_LC3_E20  <= TRANSPORT a_EQ709  ;
xor2_4825: a_EQ709 <=  n_5601  XOR n_5613;
or3_4826: n_5601 <=  n_5602  OR n_5606  OR n_5610;
and3_4827: n_5602 <=  n_5603  AND n_5604  AND n_5605;
inv_4828: n_5603  <= TRANSPORT NOT a_LC3_D22  ;
inv_4829: n_5604  <= TRANSPORT NOT a_N77_aNOT  ;
delay_4830: n_5605  <= TRANSPORT dbin(2)  ;
and2_4831: n_5606 <=  n_5607  AND n_5608;
delay_4832: n_5607  <= TRANSPORT a_N77_aNOT  ;
delay_4833: n_5608  <= TRANSPORT a_SCH2ADDRREG_F10_G  ;
and2_4834: n_5610 <=  n_5611  AND n_5612;
delay_4835: n_5611  <= TRANSPORT a_LC3_D22  ;
delay_4836: n_5612  <= TRANSPORT a_SCH2ADDRREG_F10_G  ;
and1_4837: n_5613 <=  gnd;
delay_4838: a_LC4_E20  <= TRANSPORT a_EQ710  ;
xor2_4839: a_EQ710 <=  n_5616  XOR n_5628;
or3_4840: n_5616 <=  n_5617  OR n_5621  OR n_5625;
and3_4841: n_5617 <=  n_5618  AND n_5619  AND n_5620;
inv_4842: n_5618  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_4843: n_5619  <= TRANSPORT NOT a_N2529  ;
delay_4844: n_5620  <= TRANSPORT a_LC2_A9  ;
and3_4845: n_5621 <=  n_5622  AND n_5623  AND n_5624;
inv_4846: n_5622  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_4847: n_5623  <= TRANSPORT a_N2529  ;
inv_4848: n_5624  <= TRANSPORT NOT a_LC2_A9  ;
and2_4849: n_5625 <=  n_5626  AND n_5627;
delay_4850: n_5626  <= TRANSPORT a_N2560_aNOT  ;
delay_4851: n_5627  <= TRANSPORT a_LC3_E20  ;
and1_4852: n_5628 <=  gnd;
dff_4853: DFF_a8237

    PORT MAP ( D => a_EQ1005, CLK => a_SCH2ADDRREG_F10_G_aCLK, CLRN => a_SCH2ADDRREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F10_G);
inv_4854: a_SCH2ADDRREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4855: a_EQ1005 <=  n_5635  XOR n_5642;
or2_4856: n_5635 <=  n_5636  OR n_5639;
and2_4857: n_5636 <=  n_5637  AND n_5638;
inv_4858: n_5637  <= TRANSPORT NOT a_N2527  ;
delay_4859: n_5638  <= TRANSPORT a_LC4_E20  ;
and2_4860: n_5639 <=  n_5640  AND n_5641;
delay_4861: n_5640  <= TRANSPORT a_N2527  ;
delay_4862: n_5641  <= TRANSPORT a_SCH2BAROUT_F10_G  ;
and1_4863: n_5642 <=  gnd;
delay_4864: n_5643  <= TRANSPORT clk  ;
filter_4865: FILTER_a8237

    PORT MAP (IN1 => n_5643, Y => a_SCH2ADDRREG_F10_G_aCLK);
delay_4866: a_LC4_E5  <= TRANSPORT a_EQ822  ;
xor2_4867: a_EQ822 <=  n_5647  XOR n_5655;
or2_4868: n_5647 <=  n_5648  OR n_5651;
and2_4869: n_5648 <=  n_5649  AND n_5650;
inv_4870: n_5649  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_4871: n_5650  <= TRANSPORT dbin(2)  ;
and2_4872: n_5651 <=  n_5652  AND n_5653;
delay_4873: n_5652  <= TRANSPORT a_N2573_aNOT  ;
delay_4874: n_5653  <= TRANSPORT a_SH3WRDCNTREG_F10_G  ;
and1_4875: n_5655 <=  gnd;
delay_4876: a_LC3_E5  <= TRANSPORT a_EQ823  ;
xor2_4877: a_EQ823 <=  n_5658  XOR n_5670;
or3_4878: n_5658 <=  n_5659  OR n_5662  OR n_5666;
and2_4879: n_5659 <=  n_5660  AND n_5661;
delay_4880: n_5660  <= TRANSPORT a_N965  ;
delay_4881: n_5661  <= TRANSPORT a_LC4_E5  ;
and3_4882: n_5662 <=  n_5663  AND n_5664  AND n_5665;
delay_4883: n_5663  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_4884: n_5664  <= TRANSPORT NOT a_N965  ;
inv_4885: n_5665  <= TRANSPORT NOT a_N3546  ;
and3_4886: n_5666 <=  n_5667  AND n_5668  AND n_5669;
inv_4887: n_5667  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
inv_4888: n_5668  <= TRANSPORT NOT a_N965  ;
delay_4889: n_5669  <= TRANSPORT a_N3546  ;
and1_4890: n_5670 <=  gnd;
dff_4891: DFF_a8237

    PORT MAP ( D => a_EQ1151, CLK => a_SH3WRDCNTREG_F10_G_aCLK, CLRN => a_SH3WRDCNTREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SH3WRDCNTREG_F10_G);
inv_4892: a_SH3WRDCNTREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4893: a_EQ1151 <=  n_5677  XOR n_5684;
or2_4894: n_5677 <=  n_5678  OR n_5681;
and2_4895: n_5678 <=  n_5679  AND n_5680;
inv_4896: n_5679  <= TRANSPORT NOT a_N2528  ;
delay_4897: n_5680  <= TRANSPORT a_LC3_E5  ;
and2_4898: n_5681 <=  n_5682  AND n_5683;
delay_4899: n_5682  <= TRANSPORT a_N2528  ;
delay_4900: n_5683  <= TRANSPORT a_SCH3BWORDOUT_F10_G  ;
and1_4901: n_5684 <=  gnd;
delay_4902: n_5685  <= TRANSPORT clk  ;
filter_4903: FILTER_a8237

    PORT MAP (IN1 => n_5685, Y => a_SH3WRDCNTREG_F10_G_aCLK);
delay_4904: a_LC6_E9  <= TRANSPORT a_EQ734  ;
xor2_4905: a_EQ734 <=  n_5689  XOR n_5701;
or3_4906: n_5689 <=  n_5690  OR n_5694  OR n_5698;
and3_4907: n_5690 <=  n_5691  AND n_5692  AND n_5693;
inv_4908: n_5691  <= TRANSPORT NOT a_LC3_D22  ;
inv_4909: n_5692  <= TRANSPORT NOT a_N2348  ;
delay_4910: n_5693  <= TRANSPORT dbin(2)  ;
and2_4911: n_5694 <=  n_5695  AND n_5696;
delay_4912: n_5695  <= TRANSPORT a_N2348  ;
delay_4913: n_5696  <= TRANSPORT a_SCH3ADDRREG_F10_G  ;
and2_4914: n_5698 <=  n_5699  AND n_5700;
delay_4915: n_5699  <= TRANSPORT a_LC3_D22  ;
delay_4916: n_5700  <= TRANSPORT a_SCH3ADDRREG_F10_G  ;
and1_4917: n_5701 <=  gnd;
delay_4918: a_LC4_E9  <= TRANSPORT a_EQ735  ;
xor2_4919: a_EQ735 <=  n_5704  XOR n_5716;
or3_4920: n_5704 <=  n_5705  OR n_5709  OR n_5713;
and3_4921: n_5705 <=  n_5706  AND n_5707  AND n_5708;
inv_4922: n_5706  <= TRANSPORT NOT a_N965  ;
inv_4923: n_5707  <= TRANSPORT NOT a_N2529  ;
delay_4924: n_5708  <= TRANSPORT a_LC2_A9  ;
and3_4925: n_5709 <=  n_5710  AND n_5711  AND n_5712;
inv_4926: n_5710  <= TRANSPORT NOT a_N965  ;
delay_4927: n_5711  <= TRANSPORT a_N2529  ;
inv_4928: n_5712  <= TRANSPORT NOT a_LC2_A9  ;
and2_4929: n_5713 <=  n_5714  AND n_5715;
delay_4930: n_5714  <= TRANSPORT a_N965  ;
delay_4931: n_5715  <= TRANSPORT a_LC6_E9  ;
and1_4932: n_5716 <=  gnd;
dff_4933: DFF_a8237

    PORT MAP ( D => a_EQ1069, CLK => a_SCH3ADDRREG_F10_G_aCLK, CLRN => a_SCH3ADDRREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F10_G);
inv_4934: a_SCH3ADDRREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4935: a_EQ1069 <=  n_5723  XOR n_5730;
or2_4936: n_5723 <=  n_5724  OR n_5727;
and2_4937: n_5724 <=  n_5725  AND n_5726;
inv_4938: n_5725  <= TRANSPORT NOT a_N2528  ;
delay_4939: n_5726  <= TRANSPORT a_LC4_E9  ;
and2_4940: n_5727 <=  n_5728  AND n_5729;
delay_4941: n_5728  <= TRANSPORT a_N2528  ;
delay_4942: n_5729  <= TRANSPORT a_SCH3BAROUT_F10_G  ;
and1_4943: n_5730 <=  gnd;
delay_4944: n_5731  <= TRANSPORT clk  ;
filter_4945: FILTER_a8237

    PORT MAP (IN1 => n_5731, Y => a_SCH3ADDRREG_F10_G_aCLK);
delay_4946: a_LC1_E17  <= TRANSPORT a_EQ801  ;
xor2_4947: a_EQ801 <=  n_5735  XOR n_5747;
or3_4948: n_5735 <=  n_5736  OR n_5740  OR n_5744;
and3_4949: n_5736 <=  n_5737  AND n_5738  AND n_5739;
inv_4950: n_5737  <= TRANSPORT NOT a_LC3_D22  ;
inv_4951: n_5738  <= TRANSPORT NOT a_N62_aNOT  ;
delay_4952: n_5739  <= TRANSPORT dbin(2)  ;
and2_4953: n_5740 <=  n_5741  AND n_5742;
delay_4954: n_5741  <= TRANSPORT a_N62_aNOT  ;
delay_4955: n_5742  <= TRANSPORT a_SH2WRDCNTREG_F10_G  ;
and2_4956: n_5744 <=  n_5745  AND n_5746;
delay_4957: n_5745  <= TRANSPORT a_LC3_D22  ;
delay_4958: n_5746  <= TRANSPORT a_SH2WRDCNTREG_F10_G  ;
and1_4959: n_5747 <=  gnd;
delay_4960: a_LC2_E17  <= TRANSPORT a_EQ802  ;
xor2_4961: a_EQ802 <=  n_5750  XOR n_5762;
or3_4962: n_5750 <=  n_5751  OR n_5754  OR n_5758;
and2_4963: n_5751 <=  n_5752  AND n_5753;
delay_4964: n_5752  <= TRANSPORT a_N2560_aNOT  ;
delay_4965: n_5753  <= TRANSPORT a_LC1_E17  ;
and3_4966: n_5754 <=  n_5755  AND n_5756  AND n_5757;
delay_4967: n_5755  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_4968: n_5756  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_4969: n_5757  <= TRANSPORT NOT a_N3546  ;
and3_4970: n_5758 <=  n_5759  AND n_5760  AND n_5761;
inv_4971: n_5759  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
inv_4972: n_5760  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_4973: n_5761  <= TRANSPORT a_N3546  ;
and1_4974: n_5762 <=  gnd;
dff_4975: DFF_a8237

    PORT MAP ( D => a_EQ1145, CLK => a_SH2WRDCNTREG_F10_G_aCLK, CLRN => a_SH2WRDCNTREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SH2WRDCNTREG_F10_G);
inv_4976: a_SH2WRDCNTREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_4977: a_EQ1145 <=  n_5769  XOR n_5776;
or2_4978: n_5769 <=  n_5770  OR n_5773;
and2_4979: n_5770 <=  n_5771  AND n_5772;
inv_4980: n_5771  <= TRANSPORT NOT a_N2527  ;
delay_4981: n_5772  <= TRANSPORT a_LC2_E17  ;
and2_4982: n_5773 <=  n_5774  AND n_5775;
delay_4983: n_5774  <= TRANSPORT a_N2527  ;
delay_4984: n_5775  <= TRANSPORT a_SCH2BWORDOUT_F10_G  ;
and1_4985: n_5776 <=  gnd;
delay_4986: n_5777  <= TRANSPORT clk  ;
filter_4987: FILTER_a8237

    PORT MAP (IN1 => n_5777, Y => a_SH2WRDCNTREG_F10_G_aCLK);
delay_4988: a_N2550  <= TRANSPORT a_EQ607  ;
xor2_4989: a_EQ607 <=  n_5781  XOR n_5793;
or3_4990: n_5781 <=  n_5782  OR n_5786  OR n_5790;
and3_4991: n_5782 <=  n_5783  AND n_5784  AND n_5785;
inv_4992: n_5783  <= TRANSPORT NOT a_N2529  ;
delay_4993: n_5784  <= TRANSPORT a_N2530_aNOT  ;
delay_4994: n_5785  <= TRANSPORT a_LC2_A9  ;
and3_4995: n_5786 <=  n_5787  AND n_5788  AND n_5789;
delay_4996: n_5787  <= TRANSPORT a_N2529  ;
delay_4997: n_5788  <= TRANSPORT a_N2530_aNOT  ;
inv_4998: n_5789  <= TRANSPORT NOT a_LC2_A9  ;
and2_4999: n_5790 <=  n_5791  AND n_5792;
inv_5000: n_5791  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_5001: n_5792  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and1_5002: n_5793 <=  gnd;
delay_5003: a_LC4_E11  <= TRANSPORT a_EQ681  ;
xor2_5004: a_EQ681 <=  n_5796  XOR n_5808;
or3_5005: n_5796 <=  n_5797  OR n_5801  OR n_5805;
and3_5006: n_5797 <=  n_5798  AND n_5799  AND n_5800;
inv_5007: n_5798  <= TRANSPORT NOT a_LC3_D22  ;
inv_5008: n_5799  <= TRANSPORT NOT a_N2352  ;
delay_5009: n_5800  <= TRANSPORT dbin(2)  ;
and2_5010: n_5801 <=  n_5802  AND n_5803;
delay_5011: n_5802  <= TRANSPORT a_N2352  ;
delay_5012: n_5803  <= TRANSPORT a_SCH1ADDRREG_F10_G  ;
and2_5013: n_5805 <=  n_5806  AND n_5807;
delay_5014: n_5806  <= TRANSPORT a_LC3_D22  ;
delay_5015: n_5807  <= TRANSPORT a_SCH1ADDRREG_F10_G  ;
and1_5016: n_5808 <=  gnd;
delay_5017: a_LC5_E11  <= TRANSPORT a_EQ682  ;
xor2_5018: a_EQ682 <=  n_5811  XOR n_5818;
or2_5019: n_5811 <=  n_5812  OR n_5815;
and2_5020: n_5812 <=  n_5813  AND n_5814;
inv_5021: n_5813  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_5022: n_5814  <= TRANSPORT a_N2550  ;
and2_5023: n_5815 <=  n_5816  AND n_5817;
delay_5024: n_5816  <= TRANSPORT a_N2559_aNOT  ;
delay_5025: n_5817  <= TRANSPORT a_LC4_E11  ;
and1_5026: n_5818 <=  gnd;
dff_5027: DFF_a8237

    PORT MAP ( D => a_EQ941, CLK => a_SCH1ADDRREG_F10_G_aCLK, CLRN => a_SCH1ADDRREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F10_G);
inv_5028: a_SCH1ADDRREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5029: a_EQ941 <=  n_5825  XOR n_5832;
or2_5030: n_5825 <=  n_5826  OR n_5829;
and2_5031: n_5826 <=  n_5827  AND n_5828;
inv_5032: n_5827  <= TRANSPORT NOT a_N2526  ;
delay_5033: n_5828  <= TRANSPORT a_LC5_E11  ;
and2_5034: n_5829 <=  n_5830  AND n_5831;
delay_5035: n_5830  <= TRANSPORT a_N2526  ;
delay_5036: n_5831  <= TRANSPORT a_SCH1BAROUT_F10_G  ;
and1_5037: n_5832 <=  gnd;
delay_5038: n_5833  <= TRANSPORT clk  ;
filter_5039: FILTER_a8237

    PORT MAP (IN1 => n_5833, Y => a_SCH1ADDRREG_F10_G_aCLK);
delay_5040: a_LC6_E17  <= TRANSPORT a_EQ222  ;
xor2_5041: a_EQ222 <=  n_5837  XOR n_5849;
or3_5042: n_5837 <=  n_5838  OR n_5842  OR n_5846;
and3_5043: n_5838 <=  n_5839  AND n_5840  AND n_5841;
inv_5044: n_5839  <= TRANSPORT NOT a_LC3_D22  ;
inv_5045: n_5840  <= TRANSPORT NOT a_N2353  ;
delay_5046: n_5841  <= TRANSPORT dbin(2)  ;
and2_5047: n_5842 <=  n_5843  AND n_5844;
delay_5048: n_5843  <= TRANSPORT a_N2353  ;
delay_5049: n_5844  <= TRANSPORT a_SH0WRDCNTREG_F10_G  ;
and2_5050: n_5846 <=  n_5847  AND n_5848;
delay_5051: n_5847  <= TRANSPORT a_LC3_D22  ;
delay_5052: n_5848  <= TRANSPORT a_SH0WRDCNTREG_F10_G  ;
and1_5053: n_5849 <=  gnd;
delay_5054: a_LC3_E17  <= TRANSPORT a_EQ221  ;
xor2_5055: a_EQ221 <=  n_5852  XOR n_5864;
or3_5056: n_5852 <=  n_5853  OR n_5856  OR n_5860;
and2_5057: n_5853 <=  n_5854  AND n_5855;
delay_5058: n_5854  <= TRANSPORT a_N2558_aNOT  ;
delay_5059: n_5855  <= TRANSPORT a_LC6_E17  ;
and3_5060: n_5856 <=  n_5857  AND n_5858  AND n_5859;
delay_5061: n_5857  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_5062: n_5858  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_5063: n_5859  <= TRANSPORT NOT a_N3546  ;
and3_5064: n_5860 <=  n_5861  AND n_5862  AND n_5863;
inv_5065: n_5861  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
inv_5066: n_5862  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5067: n_5863  <= TRANSPORT a_N3546  ;
and1_5068: n_5864 <=  gnd;
dff_5069: DFF_a8237

    PORT MAP ( D => a_EQ1133, CLK => a_SH0WRDCNTREG_F10_G_aCLK, CLRN => a_SH0WRDCNTREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SH0WRDCNTREG_F10_G);
inv_5070: a_SH0WRDCNTREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5071: a_EQ1133 <=  n_5871  XOR n_5878;
or2_5072: n_5871 <=  n_5872  OR n_5875;
and2_5073: n_5872 <=  n_5873  AND n_5874;
inv_5074: n_5873  <= TRANSPORT NOT a_N2525  ;
delay_5075: n_5874  <= TRANSPORT a_LC3_E17  ;
and2_5076: n_5875 <=  n_5876  AND n_5877;
delay_5077: n_5876  <= TRANSPORT a_N2525  ;
delay_5078: n_5877  <= TRANSPORT a_SCH0BWORDOUT_F10_G  ;
and1_5079: n_5878 <=  gnd;
delay_5080: n_5879  <= TRANSPORT clk  ;
filter_5081: FILTER_a8237

    PORT MAP (IN1 => n_5879, Y => a_SH0WRDCNTREG_F10_G_aCLK);
delay_5082: a_LC4_E13  <= TRANSPORT a_EQ655  ;
xor2_5083: a_EQ655 <=  n_5883  XOR n_5895;
or3_5084: n_5883 <=  n_5884  OR n_5888  OR n_5892;
and3_5085: n_5884 <=  n_5885  AND n_5886  AND n_5887;
inv_5086: n_5885  <= TRANSPORT NOT a_LC3_D22  ;
delay_5087: n_5886  <= TRANSPORT a_N2354_aNOT  ;
delay_5088: n_5887  <= TRANSPORT dbin(2)  ;
and2_5089: n_5888 <=  n_5889  AND n_5890;
inv_5090: n_5889  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_5091: n_5890  <= TRANSPORT a_SCH0ADDRREG_F10_G  ;
and2_5092: n_5892 <=  n_5893  AND n_5894;
delay_5093: n_5893  <= TRANSPORT a_LC3_D22  ;
delay_5094: n_5894  <= TRANSPORT a_SCH0ADDRREG_F10_G  ;
and1_5095: n_5895 <=  gnd;
delay_5096: a_LC5_E13  <= TRANSPORT a_EQ656  ;
xor2_5097: a_EQ656 <=  n_5898  XOR n_5905;
or2_5098: n_5898 <=  n_5899  OR n_5902;
and2_5099: n_5899 <=  n_5900  AND n_5901;
inv_5100: n_5900  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5101: n_5901  <= TRANSPORT a_N2550  ;
and2_5102: n_5902 <=  n_5903  AND n_5904;
delay_5103: n_5903  <= TRANSPORT a_N2558_aNOT  ;
delay_5104: n_5904  <= TRANSPORT a_LC4_E13  ;
and1_5105: n_5905 <=  gnd;
dff_5106: DFF_a8237

    PORT MAP ( D => a_EQ877, CLK => a_SCH0ADDRREG_F10_G_aCLK, CLRN => a_SCH0ADDRREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F10_G);
inv_5107: a_SCH0ADDRREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5108: a_EQ877 <=  n_5912  XOR n_5919;
or2_5109: n_5912 <=  n_5913  OR n_5916;
and2_5110: n_5913 <=  n_5914  AND n_5915;
inv_5111: n_5914  <= TRANSPORT NOT a_N2525  ;
delay_5112: n_5915  <= TRANSPORT a_LC5_E13  ;
and2_5113: n_5916 <=  n_5917  AND n_5918;
delay_5114: n_5917  <= TRANSPORT a_N2525  ;
delay_5115: n_5918  <= TRANSPORT a_SCH0BAROUT_F10_G  ;
and1_5116: n_5919 <=  gnd;
delay_5117: n_5920  <= TRANSPORT clk  ;
filter_5118: FILTER_a8237

    PORT MAP (IN1 => n_5920, Y => a_SCH0ADDRREG_F10_G_aCLK);
delay_5119: a_LC3_E12  <= TRANSPORT a_EQ780  ;
xor2_5120: a_EQ780 <=  n_5924  XOR n_5933;
or2_5121: n_5924 <=  n_5925  OR n_5929;
and2_5122: n_5925 <=  n_5926  AND n_5927;
delay_5123: n_5926  <= TRANSPORT a_LC2_E12  ;
delay_5124: n_5927  <= TRANSPORT a_SH1WRDCNTREG_F10_G  ;
and2_5125: n_5929 <=  n_5930  AND n_5932;
delay_5126: n_5930  <= TRANSPORT a_SCH1BWORDOUT_F10_G  ;
delay_5127: n_5932  <= TRANSPORT a_N2526  ;
and1_5128: n_5933 <=  gnd;
delay_5129: a_LC4_E12  <= TRANSPORT a_EQ781  ;
xor2_5130: a_EQ781 <=  n_5936  XOR n_5947;
or3_5131: n_5936 <=  n_5937  OR n_5939  OR n_5943;
and1_5132: n_5937 <=  n_5938;
delay_5133: n_5938  <= TRANSPORT a_LC3_E12  ;
and3_5134: n_5939 <=  n_5940  AND n_5941  AND n_5942;
delay_5135: n_5940  <= TRANSPORT a_LC4_A13_aNOT  ;
delay_5136: n_5941  <= TRANSPORT a_N460  ;
inv_5137: n_5942  <= TRANSPORT NOT a_N3546  ;
and3_5138: n_5943 <=  n_5944  AND n_5945  AND n_5946;
inv_5139: n_5944  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
delay_5140: n_5945  <= TRANSPORT a_N460  ;
delay_5141: n_5946  <= TRANSPORT a_N3546  ;
and1_5142: n_5947 <=  gnd;
dff_5143: DFF_a8237

    PORT MAP ( D => a_EQ1139, CLK => a_SH1WRDCNTREG_F10_G_aCLK, CLRN => a_SH1WRDCNTREG_F10_G_aCLRN,
          PRN => vcc, Q => a_SH1WRDCNTREG_F10_G);
inv_5144: a_SH1WRDCNTREG_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5145: a_EQ1139 <=  n_5954  XOR n_5961;
or2_5146: n_5954 <=  n_5955  OR n_5957;
and1_5147: n_5955 <=  n_5956;
delay_5148: n_5956  <= TRANSPORT a_LC4_E12  ;
and3_5149: n_5957 <=  n_5958  AND n_5959  AND n_5960;
inv_5150: n_5958  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_5151: n_5959  <= TRANSPORT a_N2595  ;
delay_5152: n_5960  <= TRANSPORT dbin(2)  ;
and1_5153: n_5961 <=  gnd;
delay_5154: n_5962  <= TRANSPORT clk  ;
filter_5155: FILTER_a8237

    PORT MAP (IN1 => n_5962, Y => a_SH1WRDCNTREG_F10_G_aCLK);
delay_5156: a_LC3_A9  <= TRANSPORT a_EQ013  ;
xor2_5157: a_EQ013 <=  n_5966  XOR n_5980;
or4_5158: n_5966 <=  n_5967  OR n_5971  OR n_5974  OR n_5977;
and3_5159: n_5967 <=  n_5968  AND n_5969  AND n_5970;
delay_5160: n_5968  <= TRANSPORT a_LC1_F10  ;
delay_5161: n_5969  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
delay_5162: n_5970  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and2_5163: n_5971 <=  n_5972  AND n_5973;
delay_5164: n_5972  <= TRANSPORT a_N757  ;
delay_5165: n_5973  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and2_5166: n_5974 <=  n_5975  AND n_5976;
delay_5167: n_5975  <= TRANSPORT a_N757  ;
delay_5168: n_5976  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
and2_5169: n_5977 <=  n_5978  AND n_5979;
delay_5170: n_5978  <= TRANSPORT a_N757  ;
delay_5171: n_5979  <= TRANSPORT a_LC1_F10  ;
and1_5172: n_5980 <=  gnd;
delay_5173: a_LC8_A9  <= TRANSPORT a_EQ007  ;
xor2_5174: a_EQ007 <=  n_5983  XOR n_5991;
or2_5175: n_5983 <=  n_5984  OR n_5988;
and2_5176: n_5984 <=  n_5985  AND n_5986;
delay_5177: n_5985  <= TRANSPORT a_LC3_A9  ;
inv_5178: n_5986  <= TRANSPORT NOT a_SADDRESSOUT_F11_G  ;
and2_5179: n_5988 <=  n_5989  AND n_5990;
inv_5180: n_5989  <= TRANSPORT NOT a_LC3_A9  ;
delay_5181: n_5990  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and1_5182: n_5991 <=  gnd;
delay_5183: a_LC1_A16  <= TRANSPORT a_EQ707  ;
xor2_5184: a_EQ707 <=  n_5994  XOR n_6002;
or2_5185: n_5994 <=  n_5995  OR n_5998;
and2_5186: n_5995 <=  n_5996  AND n_5997;
inv_5187: n_5996  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_5188: n_5997  <= TRANSPORT dbin(3)  ;
and2_5189: n_5998 <=  n_5999  AND n_6000;
delay_5190: n_5999  <= TRANSPORT a_N2583_aNOT  ;
delay_5191: n_6000  <= TRANSPORT a_SCH2ADDRREG_F11_G  ;
and1_5192: n_6002 <=  gnd;
delay_5193: a_LC2_A16  <= TRANSPORT a_EQ708  ;
xor2_5194: a_EQ708 <=  n_6005  XOR n_6017;
or3_5195: n_6005 <=  n_6006  OR n_6010  OR n_6014;
and3_5196: n_6006 <=  n_6007  AND n_6008  AND n_6009;
inv_5197: n_6007  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_5198: n_6008  <= TRANSPORT NOT a_N2529  ;
delay_5199: n_6009  <= TRANSPORT a_LC8_A9  ;
and3_5200: n_6010 <=  n_6011  AND n_6012  AND n_6013;
inv_5201: n_6011  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_5202: n_6012  <= TRANSPORT a_N2529  ;
inv_5203: n_6013  <= TRANSPORT NOT a_LC8_A9  ;
and2_5204: n_6014 <=  n_6015  AND n_6016;
delay_5205: n_6015  <= TRANSPORT a_N2560_aNOT  ;
delay_5206: n_6016  <= TRANSPORT a_LC1_A16  ;
and1_5207: n_6017 <=  gnd;
dff_5208: DFF_a8237

    PORT MAP ( D => a_EQ1006, CLK => a_SCH2ADDRREG_F11_G_aCLK, CLRN => a_SCH2ADDRREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F11_G);
inv_5209: a_SCH2ADDRREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5210: a_EQ1006 <=  n_6024  XOR n_6031;
or2_5211: n_6024 <=  n_6025  OR n_6028;
and2_5212: n_6025 <=  n_6026  AND n_6027;
inv_5213: n_6026  <= TRANSPORT NOT a_N2527  ;
delay_5214: n_6027  <= TRANSPORT a_LC2_A16  ;
and2_5215: n_6028 <=  n_6029  AND n_6030;
delay_5216: n_6029  <= TRANSPORT a_N2527  ;
delay_5217: n_6030  <= TRANSPORT a_SCH2BAROUT_F11_G  ;
and1_5218: n_6031 <=  gnd;
delay_5219: n_6032  <= TRANSPORT clk  ;
filter_5220: FILTER_a8237

    PORT MAP (IN1 => n_6032, Y => a_SCH2ADDRREG_F11_G_aCLK);
delay_5221: a_LC5_F1  <= TRANSPORT a_EQ732  ;
xor2_5222: a_EQ732 <=  n_6036  XOR n_6048;
or3_5223: n_6036 <=  n_6037  OR n_6041  OR n_6045;
and3_5224: n_6037 <=  n_6038  AND n_6039  AND n_6040;
inv_5225: n_6038  <= TRANSPORT NOT a_LC3_D22  ;
inv_5226: n_6039  <= TRANSPORT NOT a_N2348  ;
delay_5227: n_6040  <= TRANSPORT dbin(3)  ;
and2_5228: n_6041 <=  n_6042  AND n_6043;
delay_5229: n_6042  <= TRANSPORT a_N2348  ;
delay_5230: n_6043  <= TRANSPORT a_SCH3ADDRREG_F11_G  ;
and2_5231: n_6045 <=  n_6046  AND n_6047;
delay_5232: n_6046  <= TRANSPORT a_LC3_D22  ;
delay_5233: n_6047  <= TRANSPORT a_SCH3ADDRREG_F11_G  ;
and1_5234: n_6048 <=  gnd;
delay_5235: a_LC2_F1  <= TRANSPORT a_EQ733  ;
xor2_5236: a_EQ733 <=  n_6051  XOR n_6063;
or3_5237: n_6051 <=  n_6052  OR n_6056  OR n_6060;
and3_5238: n_6052 <=  n_6053  AND n_6054  AND n_6055;
inv_5239: n_6053  <= TRANSPORT NOT a_N965  ;
inv_5240: n_6054  <= TRANSPORT NOT a_N2529  ;
delay_5241: n_6055  <= TRANSPORT a_LC8_A9  ;
and3_5242: n_6056 <=  n_6057  AND n_6058  AND n_6059;
inv_5243: n_6057  <= TRANSPORT NOT a_N965  ;
delay_5244: n_6058  <= TRANSPORT a_N2529  ;
inv_5245: n_6059  <= TRANSPORT NOT a_LC8_A9  ;
and2_5246: n_6060 <=  n_6061  AND n_6062;
delay_5247: n_6061  <= TRANSPORT a_N965  ;
delay_5248: n_6062  <= TRANSPORT a_LC5_F1  ;
and1_5249: n_6063 <=  gnd;
dff_5250: DFF_a8237

    PORT MAP ( D => a_EQ1070, CLK => a_SCH3ADDRREG_F11_G_aCLK, CLRN => a_SCH3ADDRREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F11_G);
inv_5251: a_SCH3ADDRREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5252: a_EQ1070 <=  n_6070  XOR n_6077;
or2_5253: n_6070 <=  n_6071  OR n_6074;
and2_5254: n_6071 <=  n_6072  AND n_6073;
inv_5255: n_6072  <= TRANSPORT NOT a_N2528  ;
delay_5256: n_6073  <= TRANSPORT a_LC2_F1  ;
and2_5257: n_6074 <=  n_6075  AND n_6076;
delay_5258: n_6075  <= TRANSPORT a_N2528  ;
delay_5259: n_6076  <= TRANSPORT a_SCH3BAROUT_F11_G  ;
and1_5260: n_6077 <=  gnd;
delay_5261: n_6078  <= TRANSPORT clk  ;
filter_5262: FILTER_a8237

    PORT MAP (IN1 => n_6078, Y => a_SCH3ADDRREG_F11_G_aCLK);
delay_5263: a_N2551  <= TRANSPORT a_EQ608  ;
xor2_5264: a_EQ608 <=  n_6082  XOR n_6104;
or5_5265: n_6082 <=  n_6083  OR n_6087  OR n_6091  OR n_6094  OR n_6099;
and3_5266: n_6083 <=  n_6084  AND n_6085  AND n_6086;
delay_5267: n_6084  <= TRANSPORT a_N2529  ;
delay_5268: n_6085  <= TRANSPORT a_LC3_A9  ;
delay_5269: n_6086  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and3_5270: n_6087 <=  n_6088  AND n_6089  AND n_6090;
inv_5271: n_6088  <= TRANSPORT NOT a_N2529  ;
inv_5272: n_6089  <= TRANSPORT NOT a_LC3_A9  ;
delay_5273: n_6090  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and2_5274: n_6091 <=  n_6092  AND n_6093;
inv_5275: n_6092  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_5276: n_6093  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and4_5277: n_6094 <=  n_6095  AND n_6096  AND n_6097  AND n_6098;
inv_5278: n_6095  <= TRANSPORT NOT a_N2529  ;
delay_5279: n_6096  <= TRANSPORT a_N2530_aNOT  ;
delay_5280: n_6097  <= TRANSPORT a_LC3_A9  ;
inv_5281: n_6098  <= TRANSPORT NOT a_SADDRESSOUT_F11_G  ;
and4_5282: n_6099 <=  n_6100  AND n_6101  AND n_6102  AND n_6103;
delay_5283: n_6100  <= TRANSPORT a_N2529  ;
delay_5284: n_6101  <= TRANSPORT a_N2530_aNOT  ;
inv_5285: n_6102  <= TRANSPORT NOT a_LC3_A9  ;
inv_5286: n_6103  <= TRANSPORT NOT a_SADDRESSOUT_F11_G  ;
and1_5287: n_6104 <=  gnd;
delay_5288: a_LC4_A24  <= TRANSPORT a_EQ653  ;
xor2_5289: a_EQ653 <=  n_6107  XOR n_6119;
or3_5290: n_6107 <=  n_6108  OR n_6112  OR n_6116;
and3_5291: n_6108 <=  n_6109  AND n_6110  AND n_6111;
inv_5292: n_6109  <= TRANSPORT NOT a_LC3_D22  ;
delay_5293: n_6110  <= TRANSPORT a_N2354_aNOT  ;
delay_5294: n_6111  <= TRANSPORT dbin(3)  ;
and2_5295: n_6112 <=  n_6113  AND n_6114;
inv_5296: n_6113  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_5297: n_6114  <= TRANSPORT a_SCH0ADDRREG_F11_G  ;
and2_5298: n_6116 <=  n_6117  AND n_6118;
delay_5299: n_6117  <= TRANSPORT a_LC3_D22  ;
delay_5300: n_6118  <= TRANSPORT a_SCH0ADDRREG_F11_G  ;
and1_5301: n_6119 <=  gnd;
delay_5302: a_LC6_A24  <= TRANSPORT a_EQ654  ;
xor2_5303: a_EQ654 <=  n_6122  XOR n_6129;
or2_5304: n_6122 <=  n_6123  OR n_6126;
and2_5305: n_6123 <=  n_6124  AND n_6125;
inv_5306: n_6124  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5307: n_6125  <= TRANSPORT a_N2551  ;
and2_5308: n_6126 <=  n_6127  AND n_6128;
delay_5309: n_6127  <= TRANSPORT a_N2558_aNOT  ;
delay_5310: n_6128  <= TRANSPORT a_LC4_A24  ;
and1_5311: n_6129 <=  gnd;
dff_5312: DFF_a8237

    PORT MAP ( D => a_EQ878, CLK => a_SCH0ADDRREG_F11_G_aCLK, CLRN => a_SCH0ADDRREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F11_G);
inv_5313: a_SCH0ADDRREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5314: a_EQ878 <=  n_6136  XOR n_6143;
or2_5315: n_6136 <=  n_6137  OR n_6140;
and2_5316: n_6137 <=  n_6138  AND n_6139;
inv_5317: n_6138  <= TRANSPORT NOT a_N2525  ;
delay_5318: n_6139  <= TRANSPORT a_LC6_A24  ;
and2_5319: n_6140 <=  n_6141  AND n_6142;
delay_5320: n_6141  <= TRANSPORT a_N2525  ;
delay_5321: n_6142  <= TRANSPORT a_SCH0BAROUT_F11_G  ;
and1_5322: n_6143 <=  gnd;
delay_5323: n_6144  <= TRANSPORT clk  ;
filter_5324: FILTER_a8237

    PORT MAP (IN1 => n_6144, Y => a_SCH0ADDRREG_F11_G_aCLK);
delay_5325: a_LC1_A23  <= TRANSPORT a_EQ679  ;
xor2_5326: a_EQ679 <=  n_6148  XOR n_6160;
or3_5327: n_6148 <=  n_6149  OR n_6153  OR n_6157;
and3_5328: n_6149 <=  n_6150  AND n_6151  AND n_6152;
inv_5329: n_6150  <= TRANSPORT NOT a_LC3_D22  ;
inv_5330: n_6151  <= TRANSPORT NOT a_N2352  ;
delay_5331: n_6152  <= TRANSPORT dbin(3)  ;
and2_5332: n_6153 <=  n_6154  AND n_6155;
delay_5333: n_6154  <= TRANSPORT a_N2352  ;
delay_5334: n_6155  <= TRANSPORT a_SCH1ADDRREG_F11_G  ;
and2_5335: n_6157 <=  n_6158  AND n_6159;
delay_5336: n_6158  <= TRANSPORT a_LC3_D22  ;
delay_5337: n_6159  <= TRANSPORT a_SCH1ADDRREG_F11_G  ;
and1_5338: n_6160 <=  gnd;
delay_5339: a_LC2_A23  <= TRANSPORT a_EQ680  ;
xor2_5340: a_EQ680 <=  n_6163  XOR n_6170;
or2_5341: n_6163 <=  n_6164  OR n_6167;
and2_5342: n_6164 <=  n_6165  AND n_6166;
inv_5343: n_6165  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_5344: n_6166  <= TRANSPORT a_N2551  ;
and2_5345: n_6167 <=  n_6168  AND n_6169;
delay_5346: n_6168  <= TRANSPORT a_N2559_aNOT  ;
delay_5347: n_6169  <= TRANSPORT a_LC1_A23  ;
and1_5348: n_6170 <=  gnd;
dff_5349: DFF_a8237

    PORT MAP ( D => a_EQ942, CLK => a_SCH1ADDRREG_F11_G_aCLK, CLRN => a_SCH1ADDRREG_F11_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F11_G);
inv_5350: a_SCH1ADDRREG_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5351: a_EQ942 <=  n_6177  XOR n_6184;
or2_5352: n_6177 <=  n_6178  OR n_6181;
and2_5353: n_6178 <=  n_6179  AND n_6180;
inv_5354: n_6179  <= TRANSPORT NOT a_N2526  ;
delay_5355: n_6180  <= TRANSPORT a_LC2_A23  ;
and2_5356: n_6181 <=  n_6182  AND n_6183;
delay_5357: n_6182  <= TRANSPORT a_N2526  ;
delay_5358: n_6183  <= TRANSPORT a_SCH1BAROUT_F11_G  ;
and1_5359: n_6184 <=  gnd;
delay_5360: n_6185  <= TRANSPORT clk  ;
filter_5361: FILTER_a8237

    PORT MAP (IN1 => n_6185, Y => a_SCH1ADDRREG_F11_G_aCLK);
delay_5362: a_LC4_C20  <= TRANSPORT a_EQ830  ;
xor2_5363: a_EQ830 <=  n_6189  XOR n_6198;
or2_5364: n_6189 <=  n_6190  OR n_6194;
and3_5365: n_6190 <=  n_6191  AND n_6192  AND n_6193;
inv_5366: n_6191  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_5367: n_6192  <= TRANSPORT a_N1095  ;
delay_5368: n_6193  <= TRANSPORT dbin(3)  ;
and3_5369: n_6194 <=  n_6195  AND n_6196  AND n_6197;
delay_5370: n_6195  <= TRANSPORT a_N2572_aNOT  ;
delay_5371: n_6196  <= TRANSPORT a_N1095  ;
delay_5372: n_6197  <= TRANSPORT a_SCH3WRDCNTREG_F3_G  ;
and1_5373: n_6198 <=  gnd;
delay_5374: a_N1036_aNOT  <= TRANSPORT a_N1036_aNOT_aIN  ;
xor2_5375: a_N1036_aNOT_aIN <=  n_6201  XOR n_6205;
or1_5376: n_6201 <=  n_6202;
and2_5377: n_6202 <=  n_6203  AND n_6204;
inv_5378: n_6203  <= TRANSPORT NOT a_LC1_C21  ;
delay_5379: n_6204  <= TRANSPORT a_N1094  ;
and1_5380: n_6205 <=  gnd;
dff_5381: DFF_a8237

    PORT MAP ( D => a_EQ1116, CLK => a_SCH3WRDCNTREG_F3_G_aCLK, CLRN => a_SCH3WRDCNTREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F3_G);
inv_5382: a_SCH3WRDCNTREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5383: a_EQ1116 <=  n_6212  XOR n_6220;
or3_5384: n_6212 <=  n_6213  OR n_6215  OR n_6217;
and1_5385: n_6213 <=  n_6214;
delay_5386: n_6214  <= TRANSPORT a_LC4_C20  ;
and1_5387: n_6215 <=  n_6216;
delay_5388: n_6216  <= TRANSPORT a_N1036_aNOT  ;
and2_5389: n_6217 <=  n_6218  AND n_6219;
delay_5390: n_6218  <= TRANSPORT a_N2528  ;
delay_5391: n_6219  <= TRANSPORT a_SCH3BWORDOUT_F3_G  ;
and1_5392: n_6220 <=  gnd;
delay_5393: n_6221  <= TRANSPORT clk  ;
filter_5394: FILTER_a8237

    PORT MAP (IN1 => n_6221, Y => a_SCH3WRDCNTREG_F3_G_aCLK);
delay_5395: a_LC5_A9  <= TRANSPORT a_EQ008  ;
xor2_5396: a_EQ008 <=  n_6225  XOR n_6251;
or6_5397: n_6225 <=  n_6226  OR n_6231  OR n_6235  OR n_6239  OR n_6243  OR n_6247;
and3_5398: n_6226 <=  n_6227  AND n_6228  AND n_6229;
delay_5399: n_6227  <= TRANSPORT a_LC3_A9  ;
delay_5400: n_6228  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
inv_5401: n_6229  <= TRANSPORT NOT a_SADDRESSOUT_F12_G  ;
and3_5402: n_6231 <=  n_6232  AND n_6233  AND n_6234;
delay_5403: n_6232  <= TRANSPORT a_N757  ;
delay_5404: n_6233  <= TRANSPORT a_LC3_A9  ;
inv_5405: n_6234  <= TRANSPORT NOT a_SADDRESSOUT_F12_G  ;
and3_5406: n_6235 <=  n_6236  AND n_6237  AND n_6238;
delay_5407: n_6236  <= TRANSPORT a_N757  ;
delay_5408: n_6237  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
inv_5409: n_6238  <= TRANSPORT NOT a_SADDRESSOUT_F12_G  ;
and3_5410: n_6239 <=  n_6240  AND n_6241  AND n_6242;
inv_5411: n_6240  <= TRANSPORT NOT a_LC3_A9  ;
inv_5412: n_6241  <= TRANSPORT NOT a_SADDRESSOUT_F11_G  ;
delay_5413: n_6242  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and3_5414: n_6243 <=  n_6244  AND n_6245  AND n_6246;
inv_5415: n_6244  <= TRANSPORT NOT a_N757  ;
inv_5416: n_6245  <= TRANSPORT NOT a_SADDRESSOUT_F11_G  ;
delay_5417: n_6246  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and3_5418: n_6247 <=  n_6248  AND n_6249  AND n_6250;
inv_5419: n_6248  <= TRANSPORT NOT a_N757  ;
inv_5420: n_6249  <= TRANSPORT NOT a_LC3_A9  ;
delay_5421: n_6250  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and1_5422: n_6251 <=  gnd;
delay_5423: a_LC4_A14  <= TRANSPORT a_EQ705  ;
xor2_5424: a_EQ705 <=  n_6254  XOR n_6262;
or2_5425: n_6254 <=  n_6255  OR n_6258;
and2_5426: n_6255 <=  n_6256  AND n_6257;
inv_5427: n_6256  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_5428: n_6257  <= TRANSPORT dbin(4)  ;
and2_5429: n_6258 <=  n_6259  AND n_6260;
delay_5430: n_6259  <= TRANSPORT a_N2583_aNOT  ;
delay_5431: n_6260  <= TRANSPORT a_SCH2ADDRREG_F12_G  ;
and1_5432: n_6262 <=  gnd;
delay_5433: a_LC5_A14  <= TRANSPORT a_EQ706  ;
xor2_5434: a_EQ706 <=  n_6265  XOR n_6277;
or3_5435: n_6265 <=  n_6266  OR n_6270  OR n_6274;
and3_5436: n_6266 <=  n_6267  AND n_6268  AND n_6269;
inv_5437: n_6267  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_5438: n_6268  <= TRANSPORT NOT a_N2529  ;
delay_5439: n_6269  <= TRANSPORT a_LC5_A9  ;
and3_5440: n_6270 <=  n_6271  AND n_6272  AND n_6273;
inv_5441: n_6271  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_5442: n_6272  <= TRANSPORT a_N2529  ;
inv_5443: n_6273  <= TRANSPORT NOT a_LC5_A9  ;
and2_5444: n_6274 <=  n_6275  AND n_6276;
delay_5445: n_6275  <= TRANSPORT a_N2560_aNOT  ;
delay_5446: n_6276  <= TRANSPORT a_LC4_A14  ;
and1_5447: n_6277 <=  gnd;
dff_5448: DFF_a8237

    PORT MAP ( D => a_EQ1007, CLK => a_SCH2ADDRREG_F12_G_aCLK, CLRN => a_SCH2ADDRREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F12_G);
inv_5449: a_SCH2ADDRREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5450: a_EQ1007 <=  n_6284  XOR n_6291;
or2_5451: n_6284 <=  n_6285  OR n_6288;
and2_5452: n_6285 <=  n_6286  AND n_6287;
inv_5453: n_6286  <= TRANSPORT NOT a_N2527  ;
delay_5454: n_6287  <= TRANSPORT a_LC5_A14  ;
and2_5455: n_6288 <=  n_6289  AND n_6290;
delay_5456: n_6289  <= TRANSPORT a_N2527  ;
delay_5457: n_6290  <= TRANSPORT a_SCH2BAROUT_F12_G  ;
and1_5458: n_6291 <=  gnd;
delay_5459: n_6292  <= TRANSPORT clk  ;
filter_5460: FILTER_a8237

    PORT MAP (IN1 => n_6292, Y => a_SCH2ADDRREG_F12_G_aCLK);
delay_5461: a_N2552  <= TRANSPORT a_EQ609  ;
xor2_5462: a_EQ609 <=  n_6296  XOR n_6308;
or3_5463: n_6296 <=  n_6297  OR n_6301  OR n_6305;
and3_5464: n_6297 <=  n_6298  AND n_6299  AND n_6300;
inv_5465: n_6298  <= TRANSPORT NOT a_N2529  ;
delay_5466: n_6299  <= TRANSPORT a_N2530_aNOT  ;
delay_5467: n_6300  <= TRANSPORT a_LC5_A9  ;
and3_5468: n_6301 <=  n_6302  AND n_6303  AND n_6304;
delay_5469: n_6302  <= TRANSPORT a_N2529  ;
delay_5470: n_6303  <= TRANSPORT a_N2530_aNOT  ;
inv_5471: n_6304  <= TRANSPORT NOT a_LC5_A9  ;
and2_5472: n_6305 <=  n_6306  AND n_6307;
inv_5473: n_6306  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_5474: n_6307  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and1_5475: n_6308 <=  gnd;
delay_5476: a_N212  <= TRANSPORT a_N212_aIN  ;
xor2_5477: a_N212_aIN <=  n_6311  XOR n_6315;
or1_5478: n_6311 <=  n_6312;
and2_5479: n_6312 <=  n_6313  AND n_6314;
inv_5480: n_6313  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5481: n_6314  <= TRANSPORT a_N2552  ;
and1_5482: n_6315 <=  gnd;
delay_5483: a_N217  <= TRANSPORT a_EQ213  ;
xor2_5484: a_EQ213 <=  n_6318  XOR n_6328;
or2_5485: n_6318 <=  n_6319  OR n_6323;
and3_5486: n_6319 <=  n_6320  AND n_6321  AND n_6322;
inv_5487: n_6320  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_5488: n_6321  <= TRANSPORT a_N2558_aNOT  ;
delay_5489: n_6322  <= TRANSPORT dbin(4)  ;
and3_5490: n_6323 <=  n_6324  AND n_6325  AND n_6326;
delay_5491: n_6324  <= TRANSPORT a_N2587_aNOT  ;
delay_5492: n_6325  <= TRANSPORT a_N2558_aNOT  ;
delay_5493: n_6326  <= TRANSPORT a_SCH0ADDRREG_F12_G  ;
and1_5494: n_6328 <=  gnd;
dff_5495: DFF_a8237

    PORT MAP ( D => a_EQ879, CLK => a_SCH0ADDRREG_F12_G_aCLK, CLRN => a_SCH0ADDRREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F12_G);
inv_5496: a_SCH0ADDRREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5497: a_EQ879 <=  n_6335  XOR n_6345;
or3_5498: n_6335 <=  n_6336  OR n_6339  OR n_6342;
and2_5499: n_6336 <=  n_6337  AND n_6338;
inv_5500: n_6337  <= TRANSPORT NOT a_N2525  ;
delay_5501: n_6338  <= TRANSPORT a_N212  ;
and2_5502: n_6339 <=  n_6340  AND n_6341;
inv_5503: n_6340  <= TRANSPORT NOT a_N2525  ;
delay_5504: n_6341  <= TRANSPORT a_N217  ;
and2_5505: n_6342 <=  n_6343  AND n_6344;
delay_5506: n_6343  <= TRANSPORT a_N2525  ;
delay_5507: n_6344  <= TRANSPORT a_SCH0BAROUT_F12_G  ;
and1_5508: n_6345 <=  gnd;
delay_5509: n_6346  <= TRANSPORT clk  ;
filter_5510: FILTER_a8237

    PORT MAP (IN1 => n_6346, Y => a_SCH0ADDRREG_F12_G_aCLK);
delay_5511: a_LC2_A15  <= TRANSPORT a_EQ730  ;
xor2_5512: a_EQ730 <=  n_6350  XOR n_6362;
or3_5513: n_6350 <=  n_6351  OR n_6355  OR n_6359;
and3_5514: n_6351 <=  n_6352  AND n_6353  AND n_6354;
inv_5515: n_6352  <= TRANSPORT NOT a_LC3_D22  ;
inv_5516: n_6353  <= TRANSPORT NOT a_N2348  ;
delay_5517: n_6354  <= TRANSPORT dbin(4)  ;
and2_5518: n_6355 <=  n_6356  AND n_6357;
delay_5519: n_6356  <= TRANSPORT a_N2348  ;
delay_5520: n_6357  <= TRANSPORT a_SCH3ADDRREG_F12_G  ;
and2_5521: n_6359 <=  n_6360  AND n_6361;
delay_5522: n_6360  <= TRANSPORT a_LC3_D22  ;
delay_5523: n_6361  <= TRANSPORT a_SCH3ADDRREG_F12_G  ;
and1_5524: n_6362 <=  gnd;
delay_5525: a_LC1_A15  <= TRANSPORT a_EQ731  ;
xor2_5526: a_EQ731 <=  n_6365  XOR n_6377;
or3_5527: n_6365 <=  n_6366  OR n_6370  OR n_6374;
and3_5528: n_6366 <=  n_6367  AND n_6368  AND n_6369;
inv_5529: n_6367  <= TRANSPORT NOT a_N965  ;
inv_5530: n_6368  <= TRANSPORT NOT a_N2529  ;
delay_5531: n_6369  <= TRANSPORT a_LC5_A9  ;
and3_5532: n_6370 <=  n_6371  AND n_6372  AND n_6373;
inv_5533: n_6371  <= TRANSPORT NOT a_N965  ;
delay_5534: n_6372  <= TRANSPORT a_N2529  ;
inv_5535: n_6373  <= TRANSPORT NOT a_LC5_A9  ;
and2_5536: n_6374 <=  n_6375  AND n_6376;
delay_5537: n_6375  <= TRANSPORT a_N965  ;
delay_5538: n_6376  <= TRANSPORT a_LC2_A15  ;
and1_5539: n_6377 <=  gnd;
dff_5540: DFF_a8237

    PORT MAP ( D => a_EQ1071, CLK => a_SCH3ADDRREG_F12_G_aCLK, CLRN => a_SCH3ADDRREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F12_G);
inv_5541: a_SCH3ADDRREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5542: a_EQ1071 <=  n_6384  XOR n_6391;
or2_5543: n_6384 <=  n_6385  OR n_6388;
and2_5544: n_6385 <=  n_6386  AND n_6387;
inv_5545: n_6386  <= TRANSPORT NOT a_N2528  ;
delay_5546: n_6387  <= TRANSPORT a_LC1_A15  ;
and2_5547: n_6388 <=  n_6389  AND n_6390;
delay_5548: n_6389  <= TRANSPORT a_N2528  ;
delay_5549: n_6390  <= TRANSPORT a_SCH3BAROUT_F12_G  ;
and1_5550: n_6391 <=  gnd;
delay_5551: n_6392  <= TRANSPORT clk  ;
filter_5552: FILTER_a8237

    PORT MAP (IN1 => n_6392, Y => a_SCH3ADDRREG_F12_G_aCLK);
delay_5553: a_LC3_F18  <= TRANSPORT a_LC3_F18_aIN  ;
xor2_5554: a_LC3_F18_aIN <=  n_6396  XOR n_6401;
or1_5555: n_6396 <=  n_6397;
and3_5556: n_6397 <=  n_6398  AND n_6399  AND n_6400;
delay_5557: n_6398  <= TRANSPORT a_N2585_aNOT  ;
delay_5558: n_6399  <= TRANSPORT a_N2559_aNOT  ;
inv_5559: n_6400  <= TRANSPORT NOT a_N2526  ;
and1_5560: n_6401 <=  gnd;
delay_5561: a_LC8_A12  <= TRANSPORT a_EQ678  ;
xor2_5562: a_EQ678 <=  n_6404  XOR n_6412;
or2_5563: n_6404 <=  n_6405  OR n_6409;
and2_5564: n_6405 <=  n_6406  AND n_6407;
delay_5565: n_6406  <= TRANSPORT a_LC3_F18  ;
delay_5566: n_6407  <= TRANSPORT a_SCH1ADDRREG_F12_G  ;
and2_5567: n_6409 <=  n_6410  AND n_6411;
delay_5568: n_6410  <= TRANSPORT a_SCH1BAROUT_F12_G  ;
delay_5569: n_6411  <= TRANSPORT a_N2526  ;
and1_5570: n_6412 <=  gnd;
delay_5571: a_N443  <= TRANSPORT a_N443_aIN  ;
xor2_5572: a_N443_aIN <=  n_6415  XOR n_6421;
or1_5573: n_6415 <=  n_6416;
and4_5574: n_6416 <=  n_6417  AND n_6418  AND n_6419  AND n_6420;
inv_5575: n_6417  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_5576: n_6418  <= TRANSPORT a_N2559_aNOT  ;
inv_5577: n_6419  <= TRANSPORT NOT a_N2526  ;
delay_5578: n_6420  <= TRANSPORT dbin(4)  ;
and1_5579: n_6421 <=  gnd;
dff_5580: DFF_a8237

    PORT MAP ( D => a_EQ943, CLK => a_SCH1ADDRREG_F12_G_aCLK, CLRN => a_SCH1ADDRREG_F12_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F12_G);
inv_5581: a_SCH1ADDRREG_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5582: a_EQ943 <=  n_6428  XOR n_6436;
or3_5583: n_6428 <=  n_6429  OR n_6432  OR n_6434;
and2_5584: n_6429 <=  n_6430  AND n_6431;
delay_5585: n_6430  <= TRANSPORT a_N460  ;
delay_5586: n_6431  <= TRANSPORT a_N2552  ;
and1_5587: n_6432 <=  n_6433;
delay_5588: n_6433  <= TRANSPORT a_LC8_A12  ;
and1_5589: n_6434 <=  n_6435;
delay_5590: n_6435  <= TRANSPORT a_N443  ;
and1_5591: n_6436 <=  gnd;
delay_5592: n_6437  <= TRANSPORT clk  ;
filter_5593: FILTER_a8237

    PORT MAP (IN1 => n_6437, Y => a_SCH1ADDRREG_F12_G_aCLK);
delay_5594: a_N66  <= TRANSPORT a_N66_aIN  ;
xor2_5595: a_N66_aIN <=  n_6441  XOR n_6447;
or1_5596: n_6441 <=  n_6442;
and4_5597: n_6442 <=  n_6443  AND n_6444  AND n_6445  AND n_6446;
delay_5598: n_6443  <= TRANSPORT ain(3)  ;
inv_5599: n_6444  <= TRANSPORT NOT ain(2)  ;
delay_5600: n_6445  <= TRANSPORT ain(1)  ;
delay_5601: n_6446  <= TRANSPORT ain(0)  ;
and1_5602: n_6447 <=  gnd;
delay_5603: a_N2569_aNOT  <= TRANSPORT a_EQ622  ;
xor2_5604: a_EQ622 <=  n_6450  XOR n_6459;
or4_5605: n_6450 <=  n_6451  OR n_6453  OR n_6455  OR n_6457;
and1_5606: n_6451 <=  n_6452;
inv_5607: n_6452  <= TRANSPORT NOT dbin(1)  ;
and1_5608: n_6453 <=  n_6454;
delay_5609: n_6454  <= TRANSPORT dbin(0)  ;
and1_5610: n_6455 <=  n_6456;
inv_5611: n_6456  <= TRANSPORT NOT a_N66  ;
and1_5612: n_6457 <=  n_6458;
delay_5613: n_6458  <= TRANSPORT a_N87  ;
and1_5614: n_6459 <=  gnd;
dff_5615: DFF_a8237

    PORT MAP ( D => a_EQ1046, CLK => a_SCH2MODEREG_F3_G_aCLK, CLRN => a_SCH2MODEREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH2MODEREG_F3_G);
inv_5616: a_SCH2MODEREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5617: a_EQ1046 <=  n_6466  XOR n_6473;
or2_5618: n_6466 <=  n_6467  OR n_6470;
and2_5619: n_6467 <=  n_6468  AND n_6469;
delay_5620: n_6468  <= TRANSPORT a_N2569_aNOT  ;
delay_5621: n_6469  <= TRANSPORT a_SCH2MODEREG_F3_G  ;
and2_5622: n_6470 <=  n_6471  AND n_6472;
inv_5623: n_6471  <= TRANSPORT NOT a_N2569_aNOT  ;
delay_5624: n_6472  <= TRANSPORT dbin(5)  ;
and1_5625: n_6473 <=  gnd;
delay_5626: n_6474  <= TRANSPORT clk  ;
filter_5627: FILTER_a8237

    PORT MAP (IN1 => n_6474, Y => a_SCH2MODEREG_F3_G_aCLK);
delay_5628: a_N2532_aNOT  <= TRANSPORT a_N2532_aNOT_aIN  ;
xor2_5629: a_N2532_aNOT_aIN <=  n_6478  XOR n_6482;
or1_5630: n_6478 <=  n_6479;
and2_5631: n_6479 <=  n_6480  AND n_6481;
inv_5632: n_6480  <= TRANSPORT NOT dbin(0)  ;
inv_5633: n_6481  <= TRANSPORT NOT dbin(1)  ;
and1_5634: n_6482 <=  gnd;
delay_5635: a_N2567  <= TRANSPORT a_N2567_aIN  ;
xor2_5636: a_N2567_aIN <=  n_6485  XOR n_6490;
or1_5637: n_6485 <=  n_6486;
and3_5638: n_6486 <=  n_6487  AND n_6488  AND n_6489;
inv_5639: n_6487  <= TRANSPORT NOT a_N87  ;
delay_5640: n_6488  <= TRANSPORT a_N66  ;
delay_5641: n_6489  <= TRANSPORT a_N2532_aNOT  ;
and1_5642: n_6490 <=  gnd;
dff_5643: DFF_a8237

    PORT MAP ( D => a_EQ918, CLK => a_SCH0MODEREG_F3_G_aCLK, CLRN => a_SCH0MODEREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH0MODEREG_F3_G);
inv_5644: a_SCH0MODEREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5645: a_EQ918 <=  n_6497  XOR n_6504;
or2_5646: n_6497 <=  n_6498  OR n_6501;
and2_5647: n_6498 <=  n_6499  AND n_6500;
inv_5648: n_6499  <= TRANSPORT NOT a_N2567  ;
delay_5649: n_6500  <= TRANSPORT a_SCH0MODEREG_F3_G  ;
and2_5650: n_6501 <=  n_6502  AND n_6503;
delay_5651: n_6502  <= TRANSPORT a_N2567  ;
delay_5652: n_6503  <= TRANSPORT dbin(5)  ;
and1_5653: n_6504 <=  gnd;
delay_5654: n_6505  <= TRANSPORT clk  ;
filter_5655: FILTER_a8237

    PORT MAP (IN1 => n_6505, Y => a_SCH0MODEREG_F3_G_aCLK);
delay_5656: a_N84  <= TRANSPORT a_N84_aIN  ;
xor2_5657: a_N84_aIN <=  n_6509  XOR n_6513;
or1_5658: n_6509 <=  n_6510;
and2_5659: n_6510 <=  n_6511  AND n_6512;
delay_5660: n_6511  <= TRANSPORT dbin(0)  ;
inv_5661: n_6512  <= TRANSPORT NOT dbin(1)  ;
and1_5662: n_6513 <=  gnd;
delay_5663: a_N2568  <= TRANSPORT a_N2568_aIN  ;
xor2_5664: a_N2568_aIN <=  n_6516  XOR n_6521;
or1_5665: n_6516 <=  n_6517;
and3_5666: n_6517 <=  n_6518  AND n_6519  AND n_6520;
inv_5667: n_6518  <= TRANSPORT NOT a_N87  ;
delay_5668: n_6519  <= TRANSPORT a_N66  ;
delay_5669: n_6520  <= TRANSPORT a_N84  ;
and1_5670: n_6521 <=  gnd;
dff_5671: DFF_a8237

    PORT MAP ( D => a_EQ982, CLK => a_SCH1MODEREG_F3_G_aCLK, CLRN => a_SCH1MODEREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH1MODEREG_F3_G);
inv_5672: a_SCH1MODEREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5673: a_EQ982 <=  n_6528  XOR n_6535;
or2_5674: n_6528 <=  n_6529  OR n_6532;
and2_5675: n_6529 <=  n_6530  AND n_6531;
inv_5676: n_6530  <= TRANSPORT NOT a_N2568  ;
delay_5677: n_6531  <= TRANSPORT a_SCH1MODEREG_F3_G  ;
and2_5678: n_6532 <=  n_6533  AND n_6534;
delay_5679: n_6533  <= TRANSPORT a_N2568  ;
delay_5680: n_6534  <= TRANSPORT dbin(5)  ;
and1_5681: n_6535 <=  gnd;
delay_5682: n_6536  <= TRANSPORT clk  ;
filter_5683: FILTER_a8237

    PORT MAP (IN1 => n_6536, Y => a_SCH1MODEREG_F3_G_aCLK);
delay_5684: a_N2570_aNOT  <= TRANSPORT a_EQ623  ;
xor2_5685: a_EQ623 <=  n_6540  XOR n_6549;
or4_5686: n_6540 <=  n_6541  OR n_6543  OR n_6545  OR n_6547;
and1_5687: n_6541 <=  n_6542;
inv_5688: n_6542  <= TRANSPORT NOT a_N66  ;
and1_5689: n_6543 <=  n_6544;
delay_5690: n_6544  <= TRANSPORT a_N87  ;
and1_5691: n_6545 <=  n_6546;
inv_5692: n_6546  <= TRANSPORT NOT dbin(1)  ;
and1_5693: n_6547 <=  n_6548;
inv_5694: n_6548  <= TRANSPORT NOT dbin(0)  ;
and1_5695: n_6549 <=  gnd;
dff_5696: DFF_a8237

    PORT MAP ( D => a_EQ1110, CLK => a_SCH3MODEREG_F3_G_aCLK, CLRN => a_SCH3MODEREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH3MODEREG_F3_G);
inv_5697: a_SCH3MODEREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5698: a_EQ1110 <=  n_6556  XOR n_6563;
or2_5699: n_6556 <=  n_6557  OR n_6560;
and2_5700: n_6557 <=  n_6558  AND n_6559;
delay_5701: n_6558  <= TRANSPORT a_N2570_aNOT  ;
delay_5702: n_6559  <= TRANSPORT a_SCH3MODEREG_F3_G  ;
and2_5703: n_6560 <=  n_6561  AND n_6562;
inv_5704: n_6561  <= TRANSPORT NOT a_N2570_aNOT  ;
delay_5705: n_6562  <= TRANSPORT dbin(5)  ;
and1_5706: n_6563 <=  gnd;
delay_5707: n_6564  <= TRANSPORT clk  ;
filter_5708: FILTER_a8237

    PORT MAP (IN1 => n_6564, Y => a_SCH3MODEREG_F3_G_aCLK);
delay_5709: a_LC5_F8  <= TRANSPORT a_EQ263  ;
xor2_5710: a_EQ263 <=  n_6568  XOR n_6582;
or3_5711: n_6568 <=  n_6569  OR n_6573  OR n_6577;
and3_5712: n_6569 <=  n_6570  AND n_6571  AND n_6572;
inv_5713: n_6570  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5714: n_6571  <= TRANSPORT a_N3552  ;
delay_5715: n_6572  <= TRANSPORT a_N3551  ;
and3_5716: n_6573 <=  n_6574  AND n_6575  AND n_6576;
delay_5717: n_6574  <= TRANSPORT a_LC3_C13  ;
inv_5718: n_6575  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5719: n_6576  <= TRANSPORT a_N3551  ;
and4_5720: n_6577 <=  n_6578  AND n_6579  AND n_6580  AND n_6581;
inv_5721: n_6578  <= TRANSPORT NOT a_LC3_C13  ;
inv_5722: n_6579  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_5723: n_6580  <= TRANSPORT NOT a_N3552  ;
inv_5724: n_6581  <= TRANSPORT NOT a_N3551  ;
and1_5725: n_6582 <=  gnd;
delay_5726: a_LC6_F8  <= TRANSPORT a_EQ764  ;
xor2_5727: a_EQ764 <=  n_6585  XOR n_6594;
or2_5728: n_6585 <=  n_6586  OR n_6590;
and3_5729: n_6586 <=  n_6587  AND n_6588  AND n_6589;
inv_5730: n_6587  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_5731: n_6588  <= TRANSPORT a_N2558_aNOT  ;
delay_5732: n_6589  <= TRANSPORT dbin(5)  ;
and3_5733: n_6590 <=  n_6591  AND n_6592  AND n_6593;
delay_5734: n_6591  <= TRANSPORT a_N2578_aNOT  ;
delay_5735: n_6592  <= TRANSPORT a_N2558_aNOT  ;
delay_5736: n_6593  <= TRANSPORT a_SCH0WRDCNTREG_F5_G  ;
and1_5737: n_6594 <=  gnd;
dff_5738: DFF_a8237

    PORT MAP ( D => a_EQ926, CLK => a_SCH0WRDCNTREG_F5_G_aCLK, CLRN => a_SCH0WRDCNTREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F5_G);
inv_5739: a_SCH0WRDCNTREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5740: a_EQ926 <=  n_6601  XOR n_6611;
or3_5741: n_6601 <=  n_6602  OR n_6605  OR n_6608;
and2_5742: n_6602 <=  n_6603  AND n_6604;
delay_5743: n_6603  <= TRANSPORT a_N2525  ;
delay_5744: n_6604  <= TRANSPORT a_SCH0BWORDOUT_F5_G  ;
and2_5745: n_6605 <=  n_6606  AND n_6607;
inv_5746: n_6606  <= TRANSPORT NOT a_N2525  ;
delay_5747: n_6607  <= TRANSPORT a_LC5_F8  ;
and2_5748: n_6608 <=  n_6609  AND n_6610;
inv_5749: n_6609  <= TRANSPORT NOT a_N2525  ;
delay_5750: n_6610  <= TRANSPORT a_LC6_F8  ;
and1_5751: n_6611 <=  gnd;
delay_5752: n_6612  <= TRANSPORT clk  ;
filter_5753: FILTER_a8237

    PORT MAP (IN1 => n_6612, Y => a_SCH0WRDCNTREG_F5_G_aCLK);
delay_5754: a_LC8_F2  <= TRANSPORT a_EQ828  ;
xor2_5755: a_EQ828 <=  n_6616  XOR n_6625;
or2_5756: n_6616 <=  n_6617  OR n_6621;
and3_5757: n_6617 <=  n_6618  AND n_6619  AND n_6620;
inv_5758: n_6618  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_5759: n_6619  <= TRANSPORT a_N1095  ;
delay_5760: n_6620  <= TRANSPORT dbin(5)  ;
and3_5761: n_6621 <=  n_6622  AND n_6623  AND n_6624;
delay_5762: n_6622  <= TRANSPORT a_N2572_aNOT  ;
delay_5763: n_6623  <= TRANSPORT a_N1095  ;
delay_5764: n_6624  <= TRANSPORT a_SCH3WRDCNTREG_F5_G  ;
and1_5765: n_6625 <=  gnd;
delay_5766: a_N1061_aNOT  <= TRANSPORT a_EQ348  ;
xor2_5767: a_EQ348 <=  n_6628  XOR n_6642;
or3_5768: n_6628 <=  n_6629  OR n_6633  OR n_6637;
and3_5769: n_6629 <=  n_6630  AND n_6631  AND n_6632;
delay_5770: n_6630  <= TRANSPORT a_N1094  ;
delay_5771: n_6631  <= TRANSPORT a_N3552  ;
delay_5772: n_6632  <= TRANSPORT a_N3551  ;
and3_5773: n_6633 <=  n_6634  AND n_6635  AND n_6636;
delay_5774: n_6634  <= TRANSPORT a_LC3_C13  ;
delay_5775: n_6635  <= TRANSPORT a_N1094  ;
delay_5776: n_6636  <= TRANSPORT a_N3551  ;
and4_5777: n_6637 <=  n_6638  AND n_6639  AND n_6640  AND n_6641;
inv_5778: n_6638  <= TRANSPORT NOT a_LC3_C13  ;
delay_5779: n_6639  <= TRANSPORT a_N1094  ;
inv_5780: n_6640  <= TRANSPORT NOT a_N3552  ;
inv_5781: n_6641  <= TRANSPORT NOT a_N3551  ;
and1_5782: n_6642 <=  gnd;
dff_5783: DFF_a8237

    PORT MAP ( D => a_EQ1118, CLK => a_SCH3WRDCNTREG_F5_G_aCLK, CLRN => a_SCH3WRDCNTREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F5_G);
inv_5784: a_SCH3WRDCNTREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5785: a_EQ1118 <=  n_6649  XOR n_6657;
or3_5786: n_6649 <=  n_6650  OR n_6652  OR n_6654;
and1_5787: n_6650 <=  n_6651;
delay_5788: n_6651  <= TRANSPORT a_LC8_F2  ;
and1_5789: n_6652 <=  n_6653;
delay_5790: n_6653  <= TRANSPORT a_N1061_aNOT  ;
and2_5791: n_6654 <=  n_6655  AND n_6656;
delay_5792: n_6655  <= TRANSPORT a_N2528  ;
delay_5793: n_6656  <= TRANSPORT a_SCH3BWORDOUT_F5_G  ;
and1_5794: n_6657 <=  gnd;
delay_5795: n_6658  <= TRANSPORT clk  ;
filter_5796: FILTER_a8237

    PORT MAP (IN1 => n_6658, Y => a_SCH3WRDCNTREG_F5_G_aCLK);
delay_5797: a_LC3_F2  <= TRANSPORT a_EQ252  ;
xor2_5798: a_EQ252 <=  n_6662  XOR n_6676;
or3_5799: n_6662 <=  n_6663  OR n_6667  OR n_6671;
and3_5800: n_6663 <=  n_6664  AND n_6665  AND n_6666;
inv_5801: n_6664  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_5802: n_6665  <= TRANSPORT a_N3552  ;
delay_5803: n_6666  <= TRANSPORT a_N3551  ;
and3_5804: n_6667 <=  n_6668  AND n_6669  AND n_6670;
delay_5805: n_6668  <= TRANSPORT a_LC3_C13  ;
inv_5806: n_6669  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_5807: n_6670  <= TRANSPORT a_N3551  ;
and4_5808: n_6671 <=  n_6672  AND n_6673  AND n_6674  AND n_6675;
inv_5809: n_6672  <= TRANSPORT NOT a_LC3_C13  ;
inv_5810: n_6673  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_5811: n_6674  <= TRANSPORT NOT a_N3552  ;
inv_5812: n_6675  <= TRANSPORT NOT a_N3551  ;
and1_5813: n_6676 <=  gnd;
delay_5814: a_LC4_F2  <= TRANSPORT a_EQ787  ;
xor2_5815: a_EQ787 <=  n_6679  XOR n_6688;
or2_5816: n_6679 <=  n_6680  OR n_6684;
and3_5817: n_6680 <=  n_6681  AND n_6682  AND n_6683;
inv_5818: n_6681  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_5819: n_6682  <= TRANSPORT a_N2559_aNOT  ;
delay_5820: n_6683  <= TRANSPORT dbin(5)  ;
and3_5821: n_6684 <=  n_6685  AND n_6686  AND n_6687;
delay_5822: n_6685  <= TRANSPORT a_N2576_aNOT  ;
delay_5823: n_6686  <= TRANSPORT a_N2559_aNOT  ;
delay_5824: n_6687  <= TRANSPORT a_SCH1WRDCNTREG_F5_G  ;
and1_5825: n_6688 <=  gnd;
dff_5826: DFF_a8237

    PORT MAP ( D => a_EQ990, CLK => a_SCH1WRDCNTREG_F5_G_aCLK, CLRN => a_SCH1WRDCNTREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F5_G);
inv_5827: a_SCH1WRDCNTREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5828: a_EQ990 <=  n_6695  XOR n_6705;
or3_5829: n_6695 <=  n_6696  OR n_6699  OR n_6702;
and2_5830: n_6696 <=  n_6697  AND n_6698;
delay_5831: n_6697  <= TRANSPORT a_N2526  ;
delay_5832: n_6698  <= TRANSPORT a_SCH1BWORDOUT_F5_G  ;
and2_5833: n_6699 <=  n_6700  AND n_6701;
inv_5834: n_6700  <= TRANSPORT NOT a_N2526  ;
delay_5835: n_6701  <= TRANSPORT a_LC3_F2  ;
and2_5836: n_6702 <=  n_6703  AND n_6704;
inv_5837: n_6703  <= TRANSPORT NOT a_N2526  ;
delay_5838: n_6704  <= TRANSPORT a_LC4_F2  ;
and1_5839: n_6705 <=  gnd;
delay_5840: n_6706  <= TRANSPORT clk  ;
filter_5841: FILTER_a8237

    PORT MAP (IN1 => n_6706, Y => a_SCH1WRDCNTREG_F5_G_aCLK);
delay_5842: a_LC6_F24  <= TRANSPORT a_EQ808  ;
xor2_5843: a_EQ808 <=  n_6710  XOR n_6719;
or2_5844: n_6710 <=  n_6711  OR n_6715;
and3_5845: n_6711 <=  n_6712  AND n_6713  AND n_6714;
inv_5846: n_6712  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_5847: n_6713  <= TRANSPORT a_N756  ;
delay_5848: n_6714  <= TRANSPORT dbin(5)  ;
and3_5849: n_6715 <=  n_6716  AND n_6717  AND n_6718;
delay_5850: n_6716  <= TRANSPORT a_N2574_aNOT  ;
delay_5851: n_6717  <= TRANSPORT a_N756  ;
delay_5852: n_6718  <= TRANSPORT a_SCH2WRDCNTREG_F5_G  ;
and1_5853: n_6719 <=  gnd;
delay_5854: a_N833_aNOT  <= TRANSPORT a_EQ312  ;
xor2_5855: a_EQ312 <=  n_6722  XOR n_6736;
or3_5856: n_6722 <=  n_6723  OR n_6727  OR n_6731;
and3_5857: n_6723 <=  n_6724  AND n_6725  AND n_6726;
delay_5858: n_6724  <= TRANSPORT a_N858  ;
delay_5859: n_6725  <= TRANSPORT a_N3552  ;
delay_5860: n_6726  <= TRANSPORT a_N3551  ;
and3_5861: n_6727 <=  n_6728  AND n_6729  AND n_6730;
delay_5862: n_6728  <= TRANSPORT a_LC3_C13  ;
delay_5863: n_6729  <= TRANSPORT a_N858  ;
delay_5864: n_6730  <= TRANSPORT a_N3551  ;
and4_5865: n_6731 <=  n_6732  AND n_6733  AND n_6734  AND n_6735;
inv_5866: n_6732  <= TRANSPORT NOT a_LC3_C13  ;
delay_5867: n_6733  <= TRANSPORT a_N858  ;
inv_5868: n_6734  <= TRANSPORT NOT a_N3552  ;
inv_5869: n_6735  <= TRANSPORT NOT a_N3551  ;
and1_5870: n_6736 <=  gnd;
dff_5871: DFF_a8237

    PORT MAP ( D => a_EQ1054, CLK => a_SCH2WRDCNTREG_F5_G_aCLK, CLRN => a_SCH2WRDCNTREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F5_G);
inv_5872: a_SCH2WRDCNTREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5873: a_EQ1054 <=  n_6743  XOR n_6751;
or3_5874: n_6743 <=  n_6744  OR n_6746  OR n_6748;
and1_5875: n_6744 <=  n_6745;
delay_5876: n_6745  <= TRANSPORT a_LC6_F24  ;
and1_5877: n_6746 <=  n_6747;
delay_5878: n_6747  <= TRANSPORT a_N833_aNOT  ;
and2_5879: n_6748 <=  n_6749  AND n_6750;
delay_5880: n_6749  <= TRANSPORT a_N2527  ;
delay_5881: n_6750  <= TRANSPORT a_SCH2BWORDOUT_F5_G  ;
and1_5882: n_6751 <=  gnd;
delay_5883: n_6752  <= TRANSPORT clk  ;
filter_5884: FILTER_a8237

    PORT MAP (IN1 => n_6752, Y => a_SCH2WRDCNTREG_F5_G_aCLK);
delay_5885: a_LC1_E6  <= TRANSPORT a_EQ752  ;
xor2_5886: a_EQ752 <=  n_6756  XOR n_6768;
or3_5887: n_6756 <=  n_6757  OR n_6761  OR n_6765;
and3_5888: n_6757 <=  n_6758  AND n_6759  AND n_6760;
inv_5889: n_6758  <= TRANSPORT NOT a_LC3_D22  ;
inv_5890: n_6759  <= TRANSPORT NOT a_N2353  ;
delay_5891: n_6760  <= TRANSPORT dbin(5)  ;
and2_5892: n_6761 <=  n_6762  AND n_6763;
delay_5893: n_6762  <= TRANSPORT a_N2353  ;
delay_5894: n_6763  <= TRANSPORT a_SH0WRDCNTREG_F13_G  ;
and2_5895: n_6765 <=  n_6766  AND n_6767;
delay_5896: n_6766  <= TRANSPORT a_LC3_D22  ;
delay_5897: n_6767  <= TRANSPORT a_SH0WRDCNTREG_F13_G  ;
and1_5898: n_6768 <=  gnd;
delay_5899: a_LC2_E6  <= TRANSPORT a_EQ753  ;
xor2_5900: a_EQ753 <=  n_6771  XOR n_6783;
or3_5901: n_6771 <=  n_6772  OR n_6775  OR n_6779;
and2_5902: n_6772 <=  n_6773  AND n_6774;
delay_5903: n_6773  <= TRANSPORT a_N2558_aNOT  ;
delay_5904: n_6774  <= TRANSPORT a_LC1_E6  ;
and3_5905: n_6775 <=  n_6776  AND n_6777  AND n_6778;
delay_5906: n_6776  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_5907: n_6777  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_5908: n_6778  <= TRANSPORT NOT a_N3543  ;
and3_5909: n_6779 <=  n_6780  AND n_6781  AND n_6782;
inv_5910: n_6780  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
inv_5911: n_6781  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_5912: n_6782  <= TRANSPORT a_N3543  ;
and1_5913: n_6783 <=  gnd;
dff_5914: DFF_a8237

    PORT MAP ( D => a_EQ1136, CLK => a_SH0WRDCNTREG_F13_G_aCLK, CLRN => a_SH0WRDCNTREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SH0WRDCNTREG_F13_G);
inv_5915: a_SH0WRDCNTREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5916: a_EQ1136 <=  n_6790  XOR n_6797;
or2_5917: n_6790 <=  n_6791  OR n_6794;
and2_5918: n_6791 <=  n_6792  AND n_6793;
inv_5919: n_6792  <= TRANSPORT NOT a_N2525  ;
delay_5920: n_6793  <= TRANSPORT a_LC2_E6  ;
and2_5921: n_6794 <=  n_6795  AND n_6796;
delay_5922: n_6795  <= TRANSPORT a_N2525  ;
delay_5923: n_6796  <= TRANSPORT a_SCH0BWORDOUT_F13_G  ;
and1_5924: n_6797 <=  gnd;
delay_5925: n_6798  <= TRANSPORT clk  ;
filter_5926: FILTER_a8237

    PORT MAP (IN1 => n_6798, Y => a_SH0WRDCNTREG_F13_G_aCLK);
delay_5927: a_LC3_E25  <= TRANSPORT a_EQ816  ;
xor2_5928: a_EQ816 <=  n_6802  XOR n_6810;
or2_5929: n_6802 <=  n_6803  OR n_6806;
and2_5930: n_6803 <=  n_6804  AND n_6805;
inv_5931: n_6804  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_5932: n_6805  <= TRANSPORT dbin(5)  ;
and2_5933: n_6806 <=  n_6807  AND n_6808;
delay_5934: n_6807  <= TRANSPORT a_N2573_aNOT  ;
delay_5935: n_6808  <= TRANSPORT a_SH3WRDCNTREG_F13_G  ;
and1_5936: n_6810 <=  gnd;
delay_5937: a_LC4_E25  <= TRANSPORT a_EQ817  ;
xor2_5938: a_EQ817 <=  n_6813  XOR n_6825;
or3_5939: n_6813 <=  n_6814  OR n_6817  OR n_6821;
and2_5940: n_6814 <=  n_6815  AND n_6816;
delay_5941: n_6815  <= TRANSPORT a_N965  ;
delay_5942: n_6816  <= TRANSPORT a_LC3_E25  ;
and3_5943: n_6817 <=  n_6818  AND n_6819  AND n_6820;
delay_5944: n_6818  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_5945: n_6819  <= TRANSPORT NOT a_N965  ;
inv_5946: n_6820  <= TRANSPORT NOT a_N3543  ;
and3_5947: n_6821 <=  n_6822  AND n_6823  AND n_6824;
inv_5948: n_6822  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
inv_5949: n_6823  <= TRANSPORT NOT a_N965  ;
delay_5950: n_6824  <= TRANSPORT a_N3543  ;
and1_5951: n_6825 <=  gnd;
dff_5952: DFF_a8237

    PORT MAP ( D => a_EQ1154, CLK => a_SH3WRDCNTREG_F13_G_aCLK, CLRN => a_SH3WRDCNTREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SH3WRDCNTREG_F13_G);
inv_5953: a_SH3WRDCNTREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5954: a_EQ1154 <=  n_6832  XOR n_6839;
or2_5955: n_6832 <=  n_6833  OR n_6836;
and2_5956: n_6833 <=  n_6834  AND n_6835;
inv_5957: n_6834  <= TRANSPORT NOT a_N2528  ;
delay_5958: n_6835  <= TRANSPORT a_LC4_E25  ;
and2_5959: n_6836 <=  n_6837  AND n_6838;
delay_5960: n_6837  <= TRANSPORT a_N2528  ;
delay_5961: n_6838  <= TRANSPORT a_SCH3BWORDOUT_F13_G  ;
and1_5962: n_6839 <=  gnd;
delay_5963: n_6840  <= TRANSPORT clk  ;
filter_5964: FILTER_a8237

    PORT MAP (IN1 => n_6840, Y => a_SH3WRDCNTREG_F13_G_aCLK);
delay_5965: a_LC1_E19  <= TRANSPORT a_EQ774  ;
xor2_5966: a_EQ774 <=  n_6844  XOR n_6852;
or2_5967: n_6844 <=  n_6845  OR n_6848;
and2_5968: n_6845 <=  n_6846  AND n_6847;
inv_5969: n_6846  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_5970: n_6847  <= TRANSPORT dbin(5)  ;
and2_5971: n_6848 <=  n_6849  AND n_6850;
delay_5972: n_6849  <= TRANSPORT a_N2577_aNOT  ;
delay_5973: n_6850  <= TRANSPORT a_SH1WRDCNTREG_F13_G  ;
and1_5974: n_6852 <=  gnd;
delay_5975: a_LC4_E19  <= TRANSPORT a_EQ775  ;
xor2_5976: a_EQ775 <=  n_6855  XOR n_6867;
or3_5977: n_6855 <=  n_6856  OR n_6859  OR n_6863;
and2_5978: n_6856 <=  n_6857  AND n_6858;
delay_5979: n_6857  <= TRANSPORT a_N2559_aNOT  ;
delay_5980: n_6858  <= TRANSPORT a_LC1_E19  ;
and3_5981: n_6859 <=  n_6860  AND n_6861  AND n_6862;
delay_5982: n_6860  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_5983: n_6861  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_5984: n_6862  <= TRANSPORT NOT a_N3543  ;
and3_5985: n_6863 <=  n_6864  AND n_6865  AND n_6866;
inv_5986: n_6864  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
inv_5987: n_6865  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_5988: n_6866  <= TRANSPORT a_N3543  ;
and1_5989: n_6867 <=  gnd;
dff_5990: DFF_a8237

    PORT MAP ( D => a_EQ1142, CLK => a_SH1WRDCNTREG_F13_G_aCLK, CLRN => a_SH1WRDCNTREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SH1WRDCNTREG_F13_G);
inv_5991: a_SH1WRDCNTREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_5992: a_EQ1142 <=  n_6874  XOR n_6881;
or2_5993: n_6874 <=  n_6875  OR n_6878;
and2_5994: n_6875 <=  n_6876  AND n_6877;
inv_5995: n_6876  <= TRANSPORT NOT a_N2526  ;
delay_5996: n_6877  <= TRANSPORT a_LC4_E19  ;
and2_5997: n_6878 <=  n_6879  AND n_6880;
delay_5998: n_6879  <= TRANSPORT a_N2526  ;
delay_5999: n_6880  <= TRANSPORT a_SCH1BWORDOUT_F13_G  ;
and1_6000: n_6881 <=  gnd;
delay_6001: n_6882  <= TRANSPORT clk  ;
filter_6002: FILTER_a8237

    PORT MAP (IN1 => n_6882, Y => a_SH1WRDCNTREG_F13_G_aCLK);
delay_6003: a_LC1_A9  <= TRANSPORT a_EQ012  ;
xor2_6004: a_EQ012 <=  n_6886  XOR n_6900;
or4_6005: n_6886 <=  n_6887  OR n_6891  OR n_6894  OR n_6897;
and3_6006: n_6887 <=  n_6888  AND n_6889  AND n_6890;
delay_6007: n_6888  <= TRANSPORT a_LC3_A9  ;
delay_6008: n_6889  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
delay_6009: n_6890  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and2_6010: n_6891 <=  n_6892  AND n_6893;
delay_6011: n_6892  <= TRANSPORT a_N757  ;
delay_6012: n_6893  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and2_6013: n_6894 <=  n_6895  AND n_6896;
delay_6014: n_6895  <= TRANSPORT a_N757  ;
delay_6015: n_6896  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and2_6016: n_6897 <=  n_6898  AND n_6899;
delay_6017: n_6898  <= TRANSPORT a_N757  ;
delay_6018: n_6899  <= TRANSPORT a_LC3_A9  ;
and1_6019: n_6900 <=  gnd;
delay_6020: a_N2594_aNOT  <= TRANSPORT a_EQ644  ;
xor2_6021: a_EQ644 <=  n_6903  XOR n_6926;
or5_6022: n_6903 <=  n_6904  OR n_6909  OR n_6913  OR n_6916  OR n_6921;
and3_6023: n_6904 <=  n_6905  AND n_6906  AND n_6907;
delay_6024: n_6905  <= TRANSPORT a_N2529  ;
delay_6025: n_6906  <= TRANSPORT a_LC1_A9  ;
delay_6026: n_6907  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and3_6027: n_6909 <=  n_6910  AND n_6911  AND n_6912;
inv_6028: n_6910  <= TRANSPORT NOT a_N2529  ;
inv_6029: n_6911  <= TRANSPORT NOT a_LC1_A9  ;
delay_6030: n_6912  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and2_6031: n_6913 <=  n_6914  AND n_6915;
inv_6032: n_6914  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_6033: n_6915  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and4_6034: n_6916 <=  n_6917  AND n_6918  AND n_6919  AND n_6920;
inv_6035: n_6917  <= TRANSPORT NOT a_N2529  ;
delay_6036: n_6918  <= TRANSPORT a_N2530_aNOT  ;
delay_6037: n_6919  <= TRANSPORT a_LC1_A9  ;
inv_6038: n_6920  <= TRANSPORT NOT a_SADDRESSOUT_F13_G  ;
and4_6039: n_6921 <=  n_6922  AND n_6923  AND n_6924  AND n_6925;
delay_6040: n_6922  <= TRANSPORT a_N2529  ;
delay_6041: n_6923  <= TRANSPORT a_N2530_aNOT  ;
inv_6042: n_6924  <= TRANSPORT NOT a_LC1_A9  ;
inv_6043: n_6925  <= TRANSPORT NOT a_SADDRESSOUT_F13_G  ;
and1_6044: n_6926 <=  gnd;
delay_6045: a_LC7_F25  <= TRANSPORT a_EQ677  ;
xor2_6046: a_EQ677 <=  n_6929  XOR n_6937;
or2_6047: n_6929 <=  n_6930  OR n_6934;
and2_6048: n_6930 <=  n_6931  AND n_6932;
delay_6049: n_6931  <= TRANSPORT a_LC3_F18  ;
delay_6050: n_6932  <= TRANSPORT a_SCH1ADDRREG_F13_G  ;
and2_6051: n_6934 <=  n_6935  AND n_6936;
delay_6052: n_6935  <= TRANSPORT a_SCH1BAROUT_F13_G  ;
delay_6053: n_6936  <= TRANSPORT a_N2526  ;
and1_6054: n_6937 <=  gnd;
delay_6055: a_N436  <= TRANSPORT a_N436_aIN  ;
xor2_6056: a_N436_aIN <=  n_6940  XOR n_6946;
or1_6057: n_6940 <=  n_6941;
and4_6058: n_6941 <=  n_6942  AND n_6943  AND n_6944  AND n_6945;
inv_6059: n_6942  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_6060: n_6943  <= TRANSPORT a_N2559_aNOT  ;
inv_6061: n_6944  <= TRANSPORT NOT a_N2526  ;
delay_6062: n_6945  <= TRANSPORT dbin(5)  ;
and1_6063: n_6946 <=  gnd;
dff_6064: DFF_a8237

    PORT MAP ( D => a_EQ944, CLK => a_SCH1ADDRREG_F13_G_aCLK, CLRN => a_SCH1ADDRREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F13_G);
inv_6065: a_SCH1ADDRREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6066: a_EQ944 <=  n_6953  XOR n_6961;
or3_6067: n_6953 <=  n_6954  OR n_6957  OR n_6959;
and2_6068: n_6954 <=  n_6955  AND n_6956;
delay_6069: n_6955  <= TRANSPORT a_N460  ;
delay_6070: n_6956  <= TRANSPORT a_N2594_aNOT  ;
and1_6071: n_6957 <=  n_6958;
delay_6072: n_6958  <= TRANSPORT a_LC7_F25  ;
and1_6073: n_6959 <=  n_6960;
delay_6074: n_6960  <= TRANSPORT a_N436  ;
and1_6075: n_6961 <=  gnd;
delay_6076: n_6962  <= TRANSPORT clk  ;
filter_6077: FILTER_a8237

    PORT MAP (IN1 => n_6962, Y => a_SCH1ADDRREG_F13_G_aCLK);
delay_6078: a_LC5_E25  <= TRANSPORT a_EQ795  ;
xor2_6079: a_EQ795 <=  n_6966  XOR n_6978;
or3_6080: n_6966 <=  n_6967  OR n_6971  OR n_6975;
and3_6081: n_6967 <=  n_6968  AND n_6969  AND n_6970;
inv_6082: n_6968  <= TRANSPORT NOT a_LC3_D22  ;
inv_6083: n_6969  <= TRANSPORT NOT a_N62_aNOT  ;
delay_6084: n_6970  <= TRANSPORT dbin(5)  ;
and2_6085: n_6971 <=  n_6972  AND n_6973;
delay_6086: n_6972  <= TRANSPORT a_N62_aNOT  ;
delay_6087: n_6973  <= TRANSPORT a_SH2WRDCNTREG_F13_G  ;
and2_6088: n_6975 <=  n_6976  AND n_6977;
delay_6089: n_6976  <= TRANSPORT a_LC3_D22  ;
delay_6090: n_6977  <= TRANSPORT a_SH2WRDCNTREG_F13_G  ;
and1_6091: n_6978 <=  gnd;
delay_6092: a_LC6_E25  <= TRANSPORT a_EQ796  ;
xor2_6093: a_EQ796 <=  n_6981  XOR n_6993;
or3_6094: n_6981 <=  n_6982  OR n_6985  OR n_6989;
and2_6095: n_6982 <=  n_6983  AND n_6984;
delay_6096: n_6983  <= TRANSPORT a_N2560_aNOT  ;
delay_6097: n_6984  <= TRANSPORT a_LC5_E25  ;
and3_6098: n_6985 <=  n_6986  AND n_6987  AND n_6988;
delay_6099: n_6986  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_6100: n_6987  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_6101: n_6988  <= TRANSPORT NOT a_N3543  ;
and3_6102: n_6989 <=  n_6990  AND n_6991  AND n_6992;
inv_6103: n_6990  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
inv_6104: n_6991  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_6105: n_6992  <= TRANSPORT a_N3543  ;
and1_6106: n_6993 <=  gnd;
dff_6107: DFF_a8237

    PORT MAP ( D => a_EQ1148, CLK => a_SH2WRDCNTREG_F13_G_aCLK, CLRN => a_SH2WRDCNTREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SH2WRDCNTREG_F13_G);
inv_6108: a_SH2WRDCNTREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6109: a_EQ1148 <=  n_7000  XOR n_7007;
or2_6110: n_7000 <=  n_7001  OR n_7004;
and2_6111: n_7001 <=  n_7002  AND n_7003;
inv_6112: n_7002  <= TRANSPORT NOT a_N2527  ;
delay_6113: n_7003  <= TRANSPORT a_LC6_E25  ;
and2_6114: n_7004 <=  n_7005  AND n_7006;
delay_6115: n_7005  <= TRANSPORT a_N2527  ;
delay_6116: n_7006  <= TRANSPORT a_SCH2BWORDOUT_F13_G  ;
and1_6117: n_7007 <=  gnd;
delay_6118: n_7008  <= TRANSPORT clk  ;
filter_6119: FILTER_a8237

    PORT MAP (IN1 => n_7008, Y => a_SH2WRDCNTREG_F13_G_aCLK);
delay_6120: a_LC7_E3  <= TRANSPORT a_EQ009  ;
xor2_6121: a_EQ009 <=  n_7012  XOR n_7019;
or2_6122: n_7012 <=  n_7013  OR n_7016;
and2_6123: n_7013 <=  n_7014  AND n_7015;
delay_6124: n_7014  <= TRANSPORT a_LC1_A9  ;
inv_6125: n_7015  <= TRANSPORT NOT a_SADDRESSOUT_F13_G  ;
and2_6126: n_7016 <=  n_7017  AND n_7018;
inv_6127: n_7017  <= TRANSPORT NOT a_LC1_A9  ;
delay_6128: n_7018  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and1_6129: n_7019 <=  gnd;
delay_6130: a_LC1_E20  <= TRANSPORT a_EQ703  ;
xor2_6131: a_EQ703 <=  n_7022  XOR n_7030;
or2_6132: n_7022 <=  n_7023  OR n_7026;
and2_6133: n_7023 <=  n_7024  AND n_7025;
inv_6134: n_7024  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_6135: n_7025  <= TRANSPORT dbin(5)  ;
and2_6136: n_7026 <=  n_7027  AND n_7028;
delay_6137: n_7027  <= TRANSPORT a_N2583_aNOT  ;
delay_6138: n_7028  <= TRANSPORT a_SCH2ADDRREG_F13_G  ;
and1_6139: n_7030 <=  gnd;
delay_6140: a_LC2_E20  <= TRANSPORT a_EQ704  ;
xor2_6141: a_EQ704 <=  n_7033  XOR n_7045;
or3_6142: n_7033 <=  n_7034  OR n_7038  OR n_7042;
and3_6143: n_7034 <=  n_7035  AND n_7036  AND n_7037;
inv_6144: n_7035  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_6145: n_7036  <= TRANSPORT NOT a_N2529  ;
delay_6146: n_7037  <= TRANSPORT a_LC7_E3  ;
and3_6147: n_7038 <=  n_7039  AND n_7040  AND n_7041;
inv_6148: n_7039  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_6149: n_7040  <= TRANSPORT a_N2529  ;
inv_6150: n_7041  <= TRANSPORT NOT a_LC7_E3  ;
and2_6151: n_7042 <=  n_7043  AND n_7044;
delay_6152: n_7043  <= TRANSPORT a_N2560_aNOT  ;
delay_6153: n_7044  <= TRANSPORT a_LC1_E20  ;
and1_6154: n_7045 <=  gnd;
dff_6155: DFF_a8237

    PORT MAP ( D => a_EQ1008, CLK => a_SCH2ADDRREG_F13_G_aCLK, CLRN => a_SCH2ADDRREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F13_G);
inv_6156: a_SCH2ADDRREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6157: a_EQ1008 <=  n_7052  XOR n_7059;
or2_6158: n_7052 <=  n_7053  OR n_7056;
and2_6159: n_7053 <=  n_7054  AND n_7055;
inv_6160: n_7054  <= TRANSPORT NOT a_N2527  ;
delay_6161: n_7055  <= TRANSPORT a_LC2_E20  ;
and2_6162: n_7056 <=  n_7057  AND n_7058;
delay_6163: n_7057  <= TRANSPORT a_N2527  ;
delay_6164: n_7058  <= TRANSPORT a_SCH2BAROUT_F13_G  ;
and1_6165: n_7059 <=  gnd;
delay_6166: n_7060  <= TRANSPORT clk  ;
filter_6167: FILTER_a8237

    PORT MAP (IN1 => n_7060, Y => a_SCH2ADDRREG_F13_G_aCLK);
delay_6168: a_N218  <= TRANSPORT a_EQ214  ;
xor2_6169: a_EQ214 <=  n_7064  XOR n_7074;
or3_6170: n_7064 <=  n_7065  OR n_7068  OR n_7072;
and2_6171: n_7065 <=  n_7066  AND n_7067;
inv_6172: n_7066  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_6173: n_7067  <= TRANSPORT dbin(5)  ;
and2_6174: n_7068 <=  n_7069  AND n_7070;
delay_6175: n_7069  <= TRANSPORT a_N2587_aNOT  ;
delay_6176: n_7070  <= TRANSPORT a_SCH0ADDRREG_F13_G  ;
and1_6177: n_7072 <=  n_7073;
inv_6178: n_7073  <= TRANSPORT NOT a_N2558_aNOT  ;
and1_6179: n_7074 <=  gnd;
delay_6180: a_N216  <= TRANSPORT a_EQ212  ;
xor2_6181: a_EQ212 <=  n_7077  XOR n_7082;
or2_6182: n_7077 <=  n_7078  OR n_7080;
and1_6183: n_7078 <=  n_7079;
delay_6184: n_7079  <= TRANSPORT a_N2594_aNOT  ;
and1_6185: n_7080 <=  n_7081;
delay_6186: n_7081  <= TRANSPORT a_N2558_aNOT  ;
and1_6187: n_7082 <=  gnd;
dff_6188: DFF_a8237

    PORT MAP ( D => a_EQ880, CLK => a_SCH0ADDRREG_F13_G_aCLK, CLRN => a_SCH0ADDRREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F13_G);
inv_6189: a_SCH0ADDRREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6190: a_EQ880 <=  n_7089  XOR n_7097;
or2_6191: n_7089 <=  n_7090  OR n_7094;
and3_6192: n_7090 <=  n_7091  AND n_7092  AND n_7093;
inv_6193: n_7091  <= TRANSPORT NOT a_N2525  ;
delay_6194: n_7092  <= TRANSPORT a_N218  ;
delay_6195: n_7093  <= TRANSPORT a_N216  ;
and2_6196: n_7094 <=  n_7095  AND n_7096;
delay_6197: n_7095  <= TRANSPORT a_N2525  ;
delay_6198: n_7096  <= TRANSPORT a_SCH0BAROUT_F13_G  ;
and1_6199: n_7097 <=  gnd;
delay_6200: n_7098  <= TRANSPORT clk  ;
filter_6201: FILTER_a8237

    PORT MAP (IN1 => n_7098, Y => a_SCH0ADDRREG_F13_G_aCLK);
delay_6202: a_LC2_E9  <= TRANSPORT a_EQ728  ;
xor2_6203: a_EQ728 <=  n_7102  XOR n_7114;
or3_6204: n_7102 <=  n_7103  OR n_7107  OR n_7111;
and3_6205: n_7103 <=  n_7104  AND n_7105  AND n_7106;
inv_6206: n_7104  <= TRANSPORT NOT a_LC3_D22  ;
inv_6207: n_7105  <= TRANSPORT NOT a_N2348  ;
delay_6208: n_7106  <= TRANSPORT dbin(5)  ;
and2_6209: n_7107 <=  n_7108  AND n_7109;
delay_6210: n_7108  <= TRANSPORT a_N2348  ;
delay_6211: n_7109  <= TRANSPORT a_SCH3ADDRREG_F13_G  ;
and2_6212: n_7111 <=  n_7112  AND n_7113;
delay_6213: n_7112  <= TRANSPORT a_LC3_D22  ;
delay_6214: n_7113  <= TRANSPORT a_SCH3ADDRREG_F13_G  ;
and1_6215: n_7114 <=  gnd;
delay_6216: a_LC1_E9  <= TRANSPORT a_EQ729  ;
xor2_6217: a_EQ729 <=  n_7117  XOR n_7129;
or3_6218: n_7117 <=  n_7118  OR n_7122  OR n_7126;
and3_6219: n_7118 <=  n_7119  AND n_7120  AND n_7121;
inv_6220: n_7119  <= TRANSPORT NOT a_N965  ;
inv_6221: n_7120  <= TRANSPORT NOT a_N2529  ;
delay_6222: n_7121  <= TRANSPORT a_LC7_E3  ;
and3_6223: n_7122 <=  n_7123  AND n_7124  AND n_7125;
inv_6224: n_7123  <= TRANSPORT NOT a_N965  ;
delay_6225: n_7124  <= TRANSPORT a_N2529  ;
inv_6226: n_7125  <= TRANSPORT NOT a_LC7_E3  ;
and2_6227: n_7126 <=  n_7127  AND n_7128;
delay_6228: n_7127  <= TRANSPORT a_N965  ;
delay_6229: n_7128  <= TRANSPORT a_LC2_E9  ;
and1_6230: n_7129 <=  gnd;
dff_6231: DFF_a8237

    PORT MAP ( D => a_EQ1072, CLK => a_SCH3ADDRREG_F13_G_aCLK, CLRN => a_SCH3ADDRREG_F13_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F13_G);
inv_6232: a_SCH3ADDRREG_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6233: a_EQ1072 <=  n_7136  XOR n_7143;
or2_6234: n_7136 <=  n_7137  OR n_7140;
and2_6235: n_7137 <=  n_7138  AND n_7139;
inv_6236: n_7138  <= TRANSPORT NOT a_N2528  ;
delay_6237: n_7139  <= TRANSPORT a_LC1_E9  ;
and2_6238: n_7140 <=  n_7141  AND n_7142;
delay_6239: n_7141  <= TRANSPORT a_N2528  ;
delay_6240: n_7142  <= TRANSPORT a_SCH3BAROUT_F13_G  ;
and1_6241: n_7143 <=  gnd;
delay_6242: n_7144  <= TRANSPORT clk  ;
filter_6243: FILTER_a8237

    PORT MAP (IN1 => n_7144, Y => a_SCH3ADDRREG_F13_G_aCLK);
dff_6244: DFF_a8237

    PORT MAP ( D => a_EQ983, CLK => a_SCH1MODEREG_F4_G_aCLK, CLRN => a_SCH1MODEREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH1MODEREG_F4_G);
inv_6245: a_SCH1MODEREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6246: a_EQ983 <=  n_7153  XOR n_7160;
or2_6247: n_7153 <=  n_7154  OR n_7157;
and2_6248: n_7154 <=  n_7155  AND n_7156;
inv_6249: n_7155  <= TRANSPORT NOT a_N2568  ;
delay_6250: n_7156  <= TRANSPORT a_SCH1MODEREG_F4_G  ;
and2_6251: n_7157 <=  n_7158  AND n_7159;
delay_6252: n_7158  <= TRANSPORT a_N2568  ;
delay_6253: n_7159  <= TRANSPORT dbin(6)  ;
and1_6254: n_7160 <=  gnd;
delay_6255: n_7161  <= TRANSPORT clk  ;
filter_6256: FILTER_a8237

    PORT MAP (IN1 => n_7161, Y => a_SCH1MODEREG_F4_G_aCLK);
dff_6257: DFF_a8237

    PORT MAP ( D => a_EQ1047, CLK => a_SCH2MODEREG_F4_G_aCLK, CLRN => a_SCH2MODEREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH2MODEREG_F4_G);
inv_6258: a_SCH2MODEREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6259: a_EQ1047 <=  n_7170  XOR n_7177;
or2_6260: n_7170 <=  n_7171  OR n_7174;
and2_6261: n_7171 <=  n_7172  AND n_7173;
inv_6262: n_7172  <= TRANSPORT NOT a_N2569_aNOT  ;
delay_6263: n_7173  <= TRANSPORT dbin(6)  ;
and2_6264: n_7174 <=  n_7175  AND n_7176;
delay_6265: n_7175  <= TRANSPORT a_N2569_aNOT  ;
delay_6266: n_7176  <= TRANSPORT a_SCH2MODEREG_F4_G  ;
and1_6267: n_7177 <=  gnd;
delay_6268: n_7178  <= TRANSPORT clk  ;
filter_6269: FILTER_a8237

    PORT MAP (IN1 => n_7178, Y => a_SCH2MODEREG_F4_G_aCLK);
dff_6270: DFF_a8237

    PORT MAP ( D => a_EQ1111, CLK => a_SCH3MODEREG_F4_G_aCLK, CLRN => a_SCH3MODEREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH3MODEREG_F4_G);
inv_6271: a_SCH3MODEREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6272: a_EQ1111 <=  n_7187  XOR n_7194;
or2_6273: n_7187 <=  n_7188  OR n_7191;
and2_6274: n_7188 <=  n_7189  AND n_7190;
delay_6275: n_7189  <= TRANSPORT a_N2570_aNOT  ;
delay_6276: n_7190  <= TRANSPORT a_SCH3MODEREG_F4_G  ;
and2_6277: n_7191 <=  n_7192  AND n_7193;
inv_6278: n_7192  <= TRANSPORT NOT a_N2570_aNOT  ;
delay_6279: n_7193  <= TRANSPORT dbin(6)  ;
and1_6280: n_7194 <=  gnd;
delay_6281: n_7195  <= TRANSPORT clk  ;
filter_6282: FILTER_a8237

    PORT MAP (IN1 => n_7195, Y => a_SCH3MODEREG_F4_G_aCLK);
dff_6283: DFF_a8237

    PORT MAP ( D => a_EQ919, CLK => a_SCH0MODEREG_F4_G_aCLK, CLRN => a_SCH0MODEREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH0MODEREG_F4_G);
inv_6284: a_SCH0MODEREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6285: a_EQ919 <=  n_7204  XOR n_7211;
or2_6286: n_7204 <=  n_7205  OR n_7208;
and2_6287: n_7205 <=  n_7206  AND n_7207;
inv_6288: n_7206  <= TRANSPORT NOT a_N2567  ;
delay_6289: n_7207  <= TRANSPORT a_SCH0MODEREG_F4_G  ;
and2_6290: n_7208 <=  n_7209  AND n_7210;
delay_6291: n_7209  <= TRANSPORT a_N2567  ;
delay_6292: n_7210  <= TRANSPORT dbin(6)  ;
and1_6293: n_7211 <=  gnd;
delay_6294: n_7212  <= TRANSPORT clk  ;
filter_6295: FILTER_a8237

    PORT MAP (IN1 => n_7212, Y => a_SCH0MODEREG_F4_G_aCLK);
delay_6296: a_LC6_F12  <= TRANSPORT a_EQ011  ;
xor2_6297: a_EQ011 <=  n_7216  XOR n_7228;
or3_6298: n_7216 <=  n_7217  OR n_7220  OR n_7224;
and2_6299: n_7217 <=  n_7218  AND n_7219;
delay_6300: n_7218  <= TRANSPORT a_LC1_A9  ;
delay_6301: n_7219  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and3_6302: n_7220 <=  n_7221  AND n_7222  AND n_7223;
delay_6303: n_7221  <= TRANSPORT a_N2529  ;
delay_6304: n_7222  <= TRANSPORT a_N2530_aNOT  ;
delay_6305: n_7223  <= TRANSPORT a_LC1_A9  ;
and3_6306: n_7224 <=  n_7225  AND n_7226  AND n_7227;
delay_6307: n_7225  <= TRANSPORT a_N2529  ;
delay_6308: n_7226  <= TRANSPORT a_N2530_aNOT  ;
delay_6309: n_7227  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and1_6310: n_7228 <=  gnd;
delay_6311: a_LC1_F12  <= TRANSPORT a_EQ010  ;
xor2_6312: a_EQ010 <=  n_7231  XOR n_7239;
or2_6313: n_7231 <=  n_7232  OR n_7236;
and2_6314: n_7232 <=  n_7233  AND n_7234;
delay_6315: n_7233  <= TRANSPORT a_LC6_F12  ;
inv_6316: n_7234  <= TRANSPORT NOT a_SADDRESSOUT_F14_G  ;
and2_6317: n_7236 <=  n_7237  AND n_7238;
inv_6318: n_7237  <= TRANSPORT NOT a_LC6_F12  ;
delay_6319: n_7238  <= TRANSPORT a_SADDRESSOUT_F14_G  ;
and1_6320: n_7239 <=  gnd;
delay_6321: a_N2554  <= TRANSPORT a_EQ610  ;
xor2_6322: a_EQ610 <=  n_7242  XOR n_7254;
or3_6323: n_7242 <=  n_7243  OR n_7247  OR n_7251;
and3_6324: n_7243 <=  n_7244  AND n_7245  AND n_7246;
inv_6325: n_7244  <= TRANSPORT NOT a_N2529  ;
delay_6326: n_7245  <= TRANSPORT a_N2530_aNOT  ;
delay_6327: n_7246  <= TRANSPORT a_LC1_F12  ;
and3_6328: n_7247 <=  n_7248  AND n_7249  AND n_7250;
delay_6329: n_7248  <= TRANSPORT a_N2529  ;
delay_6330: n_7249  <= TRANSPORT a_N2530_aNOT  ;
inv_6331: n_7250  <= TRANSPORT NOT a_LC1_F12  ;
and2_6332: n_7251 <=  n_7252  AND n_7253;
inv_6333: n_7252  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_6334: n_7253  <= TRANSPORT a_SADDRESSOUT_F14_G  ;
and1_6335: n_7254 <=  gnd;
delay_6336: a_LC3_F7  <= TRANSPORT a_EQ651  ;
xor2_6337: a_EQ651 <=  n_7257  XOR n_7265;
or2_6338: n_7257 <=  n_7258  OR n_7261;
and2_6339: n_7258 <=  n_7259  AND n_7260;
inv_6340: n_7259  <= TRANSPORT NOT a_N2587_aNOT  ;
delay_6341: n_7260  <= TRANSPORT dbin(6)  ;
and2_6342: n_7261 <=  n_7262  AND n_7263;
delay_6343: n_7262  <= TRANSPORT a_N2587_aNOT  ;
delay_6344: n_7263  <= TRANSPORT a_SCH0ADDRREG_F14_G  ;
and1_6345: n_7265 <=  gnd;
delay_6346: a_LC4_F7  <= TRANSPORT a_EQ652  ;
xor2_6347: a_EQ652 <=  n_7268  XOR n_7275;
or2_6348: n_7268 <=  n_7269  OR n_7272;
and2_6349: n_7269 <=  n_7270  AND n_7271;
inv_6350: n_7270  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_6351: n_7271  <= TRANSPORT a_N2554  ;
and2_6352: n_7272 <=  n_7273  AND n_7274;
delay_6353: n_7273  <= TRANSPORT a_N2558_aNOT  ;
delay_6354: n_7274  <= TRANSPORT a_LC3_F7  ;
and1_6355: n_7275 <=  gnd;
dff_6356: DFF_a8237

    PORT MAP ( D => a_EQ881, CLK => a_SCH0ADDRREG_F14_G_aCLK, CLRN => a_SCH0ADDRREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F14_G);
inv_6357: a_SCH0ADDRREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6358: a_EQ881 <=  n_7282  XOR n_7289;
or2_6359: n_7282 <=  n_7283  OR n_7286;
and2_6360: n_7283 <=  n_7284  AND n_7285;
inv_6361: n_7284  <= TRANSPORT NOT a_N2525  ;
delay_6362: n_7285  <= TRANSPORT a_LC4_F7  ;
and2_6363: n_7286 <=  n_7287  AND n_7288;
delay_6364: n_7287  <= TRANSPORT a_N2525  ;
delay_6365: n_7288  <= TRANSPORT a_SCH0BAROUT_F14_G  ;
and1_6366: n_7289 <=  gnd;
delay_6367: n_7290  <= TRANSPORT clk  ;
filter_6368: FILTER_a8237

    PORT MAP (IN1 => n_7290, Y => a_SCH0ADDRREG_F14_G_aCLK);
delay_6369: a_LC1_F22  <= TRANSPORT a_EQ701  ;
xor2_6370: a_EQ701 <=  n_7294  XOR n_7302;
or2_6371: n_7294 <=  n_7295  OR n_7298;
and2_6372: n_7295 <=  n_7296  AND n_7297;
inv_6373: n_7296  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_6374: n_7297  <= TRANSPORT dbin(6)  ;
and2_6375: n_7298 <=  n_7299  AND n_7300;
delay_6376: n_7299  <= TRANSPORT a_N2583_aNOT  ;
delay_6377: n_7300  <= TRANSPORT a_SCH2ADDRREG_F14_G  ;
and1_6378: n_7302 <=  gnd;
delay_6379: a_LC3_F22  <= TRANSPORT a_EQ702  ;
xor2_6380: a_EQ702 <=  n_7305  XOR n_7312;
or2_6381: n_7305 <=  n_7306  OR n_7309;
and2_6382: n_7306 <=  n_7307  AND n_7308;
delay_6383: n_7307  <= TRANSPORT a_N756  ;
delay_6384: n_7308  <= TRANSPORT a_LC1_F22  ;
and2_6385: n_7309 <=  n_7310  AND n_7311;
delay_6386: n_7310  <= TRANSPORT a_SCH2BAROUT_F14_G  ;
delay_6387: n_7311  <= TRANSPORT a_N2527  ;
and1_6388: n_7312 <=  gnd;
dff_6389: DFF_a8237

    PORT MAP ( D => a_EQ1009, CLK => a_SCH2ADDRREG_F14_G_aCLK, CLRN => a_SCH2ADDRREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F14_G);
inv_6390: a_SCH2ADDRREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6391: a_EQ1009 <=  n_7319  XOR n_7330;
or3_6392: n_7319 <=  n_7320  OR n_7324  OR n_7328;
and3_6393: n_7320 <=  n_7321  AND n_7322  AND n_7323;
delay_6394: n_7321  <= TRANSPORT a_N858  ;
inv_6395: n_7322  <= TRANSPORT NOT a_N2529  ;
delay_6396: n_7323  <= TRANSPORT a_LC1_F12  ;
and3_6397: n_7324 <=  n_7325  AND n_7326  AND n_7327;
delay_6398: n_7325  <= TRANSPORT a_N858  ;
delay_6399: n_7326  <= TRANSPORT a_N2529  ;
inv_6400: n_7327  <= TRANSPORT NOT a_LC1_F12  ;
and1_6401: n_7328 <=  n_7329;
delay_6402: n_7329  <= TRANSPORT a_LC3_F22  ;
and1_6403: n_7330 <=  gnd;
delay_6404: n_7331  <= TRANSPORT clk  ;
filter_6405: FILTER_a8237

    PORT MAP (IN1 => n_7331, Y => a_SCH2ADDRREG_F14_G_aCLK);
delay_6406: a_LC8_F25  <= TRANSPORT a_EQ676  ;
xor2_6407: a_EQ676 <=  n_7335  XOR n_7343;
or2_6408: n_7335 <=  n_7336  OR n_7340;
and2_6409: n_7336 <=  n_7337  AND n_7338;
delay_6410: n_7337  <= TRANSPORT a_LC3_F18  ;
delay_6411: n_7338  <= TRANSPORT a_SCH1ADDRREG_F14_G  ;
and2_6412: n_7340 <=  n_7341  AND n_7342;
delay_6413: n_7341  <= TRANSPORT a_SCH1BAROUT_F14_G  ;
delay_6414: n_7342  <= TRANSPORT a_N2526  ;
and1_6415: n_7343 <=  gnd;
delay_6416: a_N440  <= TRANSPORT a_N440_aIN  ;
xor2_6417: a_N440_aIN <=  n_7346  XOR n_7352;
or1_6418: n_7346 <=  n_7347;
and4_6419: n_7347 <=  n_7348  AND n_7349  AND n_7350  AND n_7351;
inv_6420: n_7348  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_6421: n_7349  <= TRANSPORT a_N2559_aNOT  ;
inv_6422: n_7350  <= TRANSPORT NOT a_N2526  ;
delay_6423: n_7351  <= TRANSPORT dbin(6)  ;
and1_6424: n_7352 <=  gnd;
dff_6425: DFF_a8237

    PORT MAP ( D => a_EQ945, CLK => a_SCH1ADDRREG_F14_G_aCLK, CLRN => a_SCH1ADDRREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F14_G);
inv_6426: a_SCH1ADDRREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6427: a_EQ945 <=  n_7359  XOR n_7367;
or3_6428: n_7359 <=  n_7360  OR n_7363  OR n_7365;
and2_6429: n_7360 <=  n_7361  AND n_7362;
delay_6430: n_7361  <= TRANSPORT a_N460  ;
delay_6431: n_7362  <= TRANSPORT a_N2554  ;
and1_6432: n_7363 <=  n_7364;
delay_6433: n_7364  <= TRANSPORT a_LC8_F25  ;
and1_6434: n_7365 <=  n_7366;
delay_6435: n_7366  <= TRANSPORT a_N440  ;
and1_6436: n_7367 <=  gnd;
delay_6437: n_7368  <= TRANSPORT clk  ;
filter_6438: FILTER_a8237

    PORT MAP (IN1 => n_7368, Y => a_SCH1ADDRREG_F14_G_aCLK);
delay_6439: a_LC4_F1  <= TRANSPORT a_EQ726  ;
xor2_6440: a_EQ726 <=  n_7372  XOR n_7384;
or3_6441: n_7372 <=  n_7373  OR n_7377  OR n_7381;
and3_6442: n_7373 <=  n_7374  AND n_7375  AND n_7376;
inv_6443: n_7374  <= TRANSPORT NOT a_LC3_D22  ;
inv_6444: n_7375  <= TRANSPORT NOT a_N2348  ;
delay_6445: n_7376  <= TRANSPORT dbin(6)  ;
and2_6446: n_7377 <=  n_7378  AND n_7379;
delay_6447: n_7378  <= TRANSPORT a_N2348  ;
delay_6448: n_7379  <= TRANSPORT a_SCH3ADDRREG_F14_G  ;
and2_6449: n_7381 <=  n_7382  AND n_7383;
delay_6450: n_7382  <= TRANSPORT a_LC3_D22  ;
delay_6451: n_7383  <= TRANSPORT a_SCH3ADDRREG_F14_G  ;
and1_6452: n_7384 <=  gnd;
delay_6453: a_LC3_F1  <= TRANSPORT a_EQ727  ;
xor2_6454: a_EQ727 <=  n_7387  XOR n_7399;
or3_6455: n_7387 <=  n_7388  OR n_7392  OR n_7396;
and3_6456: n_7388 <=  n_7389  AND n_7390  AND n_7391;
inv_6457: n_7389  <= TRANSPORT NOT a_N965  ;
inv_6458: n_7390  <= TRANSPORT NOT a_N2529  ;
delay_6459: n_7391  <= TRANSPORT a_LC1_F12  ;
and3_6460: n_7392 <=  n_7393  AND n_7394  AND n_7395;
inv_6461: n_7393  <= TRANSPORT NOT a_N965  ;
delay_6462: n_7394  <= TRANSPORT a_N2529  ;
inv_6463: n_7395  <= TRANSPORT NOT a_LC1_F12  ;
and2_6464: n_7396 <=  n_7397  AND n_7398;
delay_6465: n_7397  <= TRANSPORT a_N965  ;
delay_6466: n_7398  <= TRANSPORT a_LC4_F1  ;
and1_6467: n_7399 <=  gnd;
dff_6468: DFF_a8237

    PORT MAP ( D => a_EQ1073, CLK => a_SCH3ADDRREG_F14_G_aCLK, CLRN => a_SCH3ADDRREG_F14_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F14_G);
inv_6469: a_SCH3ADDRREG_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6470: a_EQ1073 <=  n_7406  XOR n_7413;
or2_6471: n_7406 <=  n_7407  OR n_7410;
and2_6472: n_7407 <=  n_7408  AND n_7409;
inv_6473: n_7408  <= TRANSPORT NOT a_N2528  ;
delay_6474: n_7409  <= TRANSPORT a_LC3_F1  ;
and2_6475: n_7410 <=  n_7411  AND n_7412;
delay_6476: n_7411  <= TRANSPORT a_N2528  ;
delay_6477: n_7412  <= TRANSPORT a_SCH3BAROUT_F14_G  ;
and1_6478: n_7413 <=  gnd;
delay_6479: n_7414  <= TRANSPORT clk  ;
filter_6480: FILTER_a8237

    PORT MAP (IN1 => n_7414, Y => a_SCH3ADDRREG_F14_G_aCLK);
delay_6481: a_LC4_D2  <= TRANSPORT a_EQ826  ;
xor2_6482: a_EQ826 <=  n_7418  XOR n_7428;
or2_6483: n_7418 <=  n_7419  OR n_7423;
and3_6484: n_7419 <=  n_7420  AND n_7421  AND n_7422;
inv_6485: n_7420  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_6486: n_7421  <= TRANSPORT a_N1095  ;
delay_6487: n_7422  <= TRANSPORT dbin(7)  ;
and3_6488: n_7423 <=  n_7424  AND n_7425  AND n_7426;
delay_6489: n_7424  <= TRANSPORT a_N2572_aNOT  ;
delay_6490: n_7425  <= TRANSPORT a_N1095  ;
delay_6491: n_7426  <= TRANSPORT a_SCH3WRDCNTREG_F7_G  ;
and1_6492: n_7428 <=  gnd;
delay_6493: a_N1038_aNOT  <= TRANSPORT a_EQ345  ;
xor2_6494: a_EQ345 <=  n_7431  XOR n_7440;
or2_6495: n_7431 <=  n_7432  OR n_7436;
and3_6496: n_7432 <=  n_7433  AND n_7434  AND n_7435;
delay_6497: n_7433  <= TRANSPORT a_LC8_F13_aNOT  ;
delay_6498: n_7434  <= TRANSPORT a_N1094  ;
inv_6499: n_7435  <= TRANSPORT NOT a_N3549  ;
and3_6500: n_7436 <=  n_7437  AND n_7438  AND n_7439;
inv_6501: n_7437  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
delay_6502: n_7438  <= TRANSPORT a_N1094  ;
delay_6503: n_7439  <= TRANSPORT a_N3549  ;
and1_6504: n_7440 <=  gnd;
dff_6505: DFF_a8237

    PORT MAP ( D => a_EQ1120, CLK => a_SCH3WRDCNTREG_F7_G_aCLK, CLRN => a_SCH3WRDCNTREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH3WRDCNTREG_F7_G);
inv_6506: a_SCH3WRDCNTREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6507: a_EQ1120 <=  n_7447  XOR n_7455;
or3_6508: n_7447 <=  n_7448  OR n_7450  OR n_7452;
and1_6509: n_7448 <=  n_7449;
delay_6510: n_7449  <= TRANSPORT a_LC4_D2  ;
and1_6511: n_7450 <=  n_7451;
delay_6512: n_7451  <= TRANSPORT a_N1038_aNOT  ;
and2_6513: n_7452 <=  n_7453  AND n_7454;
delay_6514: n_7453  <= TRANSPORT a_N2528  ;
delay_6515: n_7454  <= TRANSPORT a_SCH3BWORDOUT_F7_G  ;
and1_6516: n_7455 <=  gnd;
delay_6517: n_7456  <= TRANSPORT clk  ;
filter_6518: FILTER_a8237

    PORT MAP (IN1 => n_7456, Y => a_SCH3WRDCNTREG_F7_G_aCLK);
delay_6519: a_N782_aNOT  <= TRANSPORT a_EQ298  ;
xor2_6520: a_EQ298 <=  n_7460  XOR n_7468;
or2_6521: n_7460 <=  n_7461  OR n_7464;
and2_6522: n_7461 <=  n_7462  AND n_7463;
inv_6523: n_7462  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_6524: n_7463  <= TRANSPORT dbin(7)  ;
and2_6525: n_7464 <=  n_7465  AND n_7466;
delay_6526: n_7465  <= TRANSPORT a_N2574_aNOT  ;
delay_6527: n_7466  <= TRANSPORT a_SCH2WRDCNTREG_F7_G  ;
and1_6528: n_7468 <=  gnd;
delay_6529: a_LC5_D5  <= TRANSPORT a_EQ806  ;
xor2_6530: a_EQ806 <=  n_7471  XOR n_7483;
or3_6531: n_7471 <=  n_7472  OR n_7475  OR n_7479;
and2_6532: n_7472 <=  n_7473  AND n_7474;
delay_6533: n_7473  <= TRANSPORT a_N2560_aNOT  ;
delay_6534: n_7474  <= TRANSPORT a_N782_aNOT  ;
and3_6535: n_7475 <=  n_7476  AND n_7477  AND n_7478;
delay_6536: n_7476  <= TRANSPORT a_LC8_F13_aNOT  ;
inv_6537: n_7477  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_6538: n_7478  <= TRANSPORT NOT a_N3549  ;
and3_6539: n_7479 <=  n_7480  AND n_7481  AND n_7482;
inv_6540: n_7480  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
inv_6541: n_7481  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_6542: n_7482  <= TRANSPORT a_N3549  ;
and1_6543: n_7483 <=  gnd;
dff_6544: DFF_a8237

    PORT MAP ( D => a_EQ1056, CLK => a_SCH2WRDCNTREG_F7_G_aCLK, CLRN => a_SCH2WRDCNTREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH2WRDCNTREG_F7_G);
inv_6545: a_SCH2WRDCNTREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6546: a_EQ1056 <=  n_7490  XOR n_7497;
or2_6547: n_7490 <=  n_7491  OR n_7494;
and2_6548: n_7491 <=  n_7492  AND n_7493;
inv_6549: n_7492  <= TRANSPORT NOT a_N2527  ;
delay_6550: n_7493  <= TRANSPORT a_LC5_D5  ;
and2_6551: n_7494 <=  n_7495  AND n_7496;
delay_6552: n_7495  <= TRANSPORT a_N2527  ;
delay_6553: n_7496  <= TRANSPORT a_SCH2BWORDOUT_F7_G  ;
and1_6554: n_7497 <=  gnd;
delay_6555: n_7498  <= TRANSPORT clk  ;
filter_6556: FILTER_a8237

    PORT MAP (IN1 => n_7498, Y => a_SCH2WRDCNTREG_F7_G_aCLK);
delay_6557: a_N646_aNOT  <= TRANSPORT a_EQ278  ;
xor2_6558: a_EQ278 <=  n_7502  XOR n_7510;
or2_6559: n_7502 <=  n_7503  OR n_7506;
and2_6560: n_7503 <=  n_7504  AND n_7505;
inv_6561: n_7504  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_6562: n_7505  <= TRANSPORT dbin(7)  ;
and2_6563: n_7506 <=  n_7507  AND n_7508;
delay_6564: n_7507  <= TRANSPORT a_N2576_aNOT  ;
delay_6565: n_7508  <= TRANSPORT a_SCH1WRDCNTREG_F7_G  ;
and1_6566: n_7510 <=  gnd;
delay_6567: a_LC4_D11  <= TRANSPORT a_EQ784  ;
xor2_6568: a_EQ784 <=  n_7513  XOR n_7521;
or2_6569: n_7513 <=  n_7514  OR n_7518;
and3_6570: n_7514 <=  n_7515  AND n_7516  AND n_7517;
delay_6571: n_7515  <= TRANSPORT a_N2559_aNOT  ;
inv_6572: n_7516  <= TRANSPORT NOT a_N2526  ;
delay_6573: n_7517  <= TRANSPORT a_N646_aNOT  ;
and2_6574: n_7518 <=  n_7519  AND n_7520;
delay_6575: n_7519  <= TRANSPORT a_SCH1BWORDOUT_F7_G  ;
delay_6576: n_7520  <= TRANSPORT a_N2526  ;
and1_6577: n_7521 <=  gnd;
dff_6578: DFF_a8237

    PORT MAP ( D => a_EQ992, CLK => a_SCH1WRDCNTREG_F7_G_aCLK, CLRN => a_SCH1WRDCNTREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH1WRDCNTREG_F7_G);
inv_6579: a_SCH1WRDCNTREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6580: a_EQ992 <=  n_7528  XOR n_7539;
or3_6581: n_7528 <=  n_7529  OR n_7531  OR n_7535;
and1_6582: n_7529 <=  n_7530;
delay_6583: n_7530  <= TRANSPORT a_LC4_D11  ;
and3_6584: n_7531 <=  n_7532  AND n_7533  AND n_7534;
delay_6585: n_7532  <= TRANSPORT a_LC8_F13_aNOT  ;
delay_6586: n_7533  <= TRANSPORT a_N460  ;
inv_6587: n_7534  <= TRANSPORT NOT a_N3549  ;
and3_6588: n_7535 <=  n_7536  AND n_7537  AND n_7538;
inv_6589: n_7536  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
delay_6590: n_7537  <= TRANSPORT a_N460  ;
delay_6591: n_7538  <= TRANSPORT a_N3549  ;
and1_6592: n_7539 <=  gnd;
delay_6593: n_7540  <= TRANSPORT clk  ;
filter_6594: FILTER_a8237

    PORT MAP (IN1 => n_7540, Y => a_SCH1WRDCNTREG_F7_G_aCLK);
delay_6595: a_LC4_D9  <= TRANSPORT a_EQ760  ;
xor2_6596: a_EQ760 <=  n_7544  XOR n_7552;
or2_6597: n_7544 <=  n_7545  OR n_7548;
and2_6598: n_7545 <=  n_7546  AND n_7547;
inv_6599: n_7546  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_6600: n_7547  <= TRANSPORT dbin(7)  ;
and2_6601: n_7548 <=  n_7549  AND n_7550;
delay_6602: n_7549  <= TRANSPORT a_N2578_aNOT  ;
delay_6603: n_7550  <= TRANSPORT a_SCH0WRDCNTREG_F7_G  ;
and1_6604: n_7552 <=  gnd;
delay_6605: a_LC5_D9  <= TRANSPORT a_EQ761  ;
xor2_6606: a_EQ761 <=  n_7555  XOR n_7567;
or3_6607: n_7555 <=  n_7556  OR n_7559  OR n_7563;
and2_6608: n_7556 <=  n_7557  AND n_7558;
delay_6609: n_7557  <= TRANSPORT a_N2558_aNOT  ;
delay_6610: n_7558  <= TRANSPORT a_LC4_D9  ;
and3_6611: n_7559 <=  n_7560  AND n_7561  AND n_7562;
delay_6612: n_7560  <= TRANSPORT a_LC8_F13_aNOT  ;
inv_6613: n_7561  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_6614: n_7562  <= TRANSPORT NOT a_N3549  ;
and3_6615: n_7563 <=  n_7564  AND n_7565  AND n_7566;
inv_6616: n_7564  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
inv_6617: n_7565  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_6618: n_7566  <= TRANSPORT a_N3549  ;
and1_6619: n_7567 <=  gnd;
dff_6620: DFF_a8237

    PORT MAP ( D => a_EQ928, CLK => a_SCH0WRDCNTREG_F7_G_aCLK, CLRN => a_SCH0WRDCNTREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH0WRDCNTREG_F7_G);
inv_6621: a_SCH0WRDCNTREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6622: a_EQ928 <=  n_7574  XOR n_7581;
or2_6623: n_7574 <=  n_7575  OR n_7578;
and2_6624: n_7575 <=  n_7576  AND n_7577;
inv_6625: n_7576  <= TRANSPORT NOT a_N2525  ;
delay_6626: n_7577  <= TRANSPORT a_LC5_D9  ;
and2_6627: n_7578 <=  n_7579  AND n_7580;
delay_6628: n_7579  <= TRANSPORT a_N2525  ;
delay_6629: n_7580  <= TRANSPORT a_SCH0BWORDOUT_F7_G  ;
and1_6630: n_7581 <=  gnd;
delay_6631: n_7582  <= TRANSPORT clk  ;
filter_6632: FILTER_a8237

    PORT MAP (IN1 => n_7582, Y => a_SCH0WRDCNTREG_F7_G_aCLK);
delay_6633: a_LC3_F12  <= TRANSPORT a_EQ834  ;
xor2_6634: a_EQ834 <=  n_7586  XOR n_7599;
or3_6635: n_7586 <=  n_7587  OR n_7591  OR n_7595;
and3_6636: n_7587 <=  n_7588  AND n_7589  AND n_7590;
delay_6637: n_7588  <= TRANSPORT a_N2529  ;
inv_6638: n_7589  <= TRANSPORT NOT a_LC1_F12  ;
inv_6639: n_7590  <= TRANSPORT NOT a_SADDRESSOUT_F14_G  ;
and3_6640: n_7591 <=  n_7592  AND n_7593  AND n_7594;
delay_6641: n_7592  <= TRANSPORT a_N2529  ;
inv_6642: n_7593  <= TRANSPORT NOT a_LC6_F12  ;
inv_6643: n_7594  <= TRANSPORT NOT a_LC1_F12  ;
and3_6644: n_7595 <=  n_7596  AND n_7597  AND n_7598;
inv_6645: n_7596  <= TRANSPORT NOT a_N2529  ;
delay_6646: n_7597  <= TRANSPORT a_LC6_F12  ;
delay_6647: n_7598  <= TRANSPORT a_SADDRESSOUT_F14_G  ;
and1_6648: n_7599 <=  gnd;
delay_6649: a_N3045  <= TRANSPORT a_EQ835  ;
xor2_6650: a_EQ835 <=  n_7602  XOR n_7610;
or2_6651: n_7602 <=  n_7603  OR n_7607;
and2_6652: n_7603 <=  n_7604  AND n_7605;
delay_6653: n_7604  <= TRANSPORT a_LC3_F12  ;
inv_6654: n_7605  <= TRANSPORT NOT a_SADDRESSOUT_F15_G  ;
and2_6655: n_7607 <=  n_7608  AND n_7609;
inv_6656: n_7608  <= TRANSPORT NOT a_LC3_F12  ;
delay_6657: n_7609  <= TRANSPORT a_SADDRESSOUT_F15_G  ;
and1_6658: n_7610 <=  gnd;
delay_6659: a_LC6_D5  <= TRANSPORT a_EQ700  ;
xor2_6660: a_EQ700 <=  n_7613  XOR n_7622;
or2_6661: n_7613 <=  n_7614  OR n_7617;
and2_6662: n_7614 <=  n_7615  AND n_7616;
inv_6663: n_7615  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_6664: n_7616  <= TRANSPORT a_N3045  ;
and3_6665: n_7617 <=  n_7618  AND n_7619  AND n_7620;
delay_6666: n_7618  <= TRANSPORT a_N2583_aNOT  ;
delay_6667: n_7619  <= TRANSPORT a_N2560_aNOT  ;
delay_6668: n_7620  <= TRANSPORT a_SCH2ADDRREG_F15_G  ;
and1_6669: n_7622 <=  gnd;
delay_6670: a_N818  <= TRANSPORT a_N818_aIN  ;
xor2_6671: a_N818_aIN <=  n_7625  XOR n_7630;
or1_6672: n_7625 <=  n_7626;
and3_6673: n_7626 <=  n_7627  AND n_7628  AND n_7629;
inv_6674: n_7627  <= TRANSPORT NOT a_N2583_aNOT  ;
delay_6675: n_7628  <= TRANSPORT a_N756  ;
delay_6676: n_7629  <= TRANSPORT dbin(7)  ;
and1_6677: n_7630 <=  gnd;
dff_6678: DFF_a8237

    PORT MAP ( D => a_EQ1010, CLK => a_SCH2ADDRREG_F15_G_aCLK, CLRN => a_SCH2ADDRREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F15_G);
inv_6679: a_SCH2ADDRREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6680: a_EQ1010 <=  n_7637  XOR n_7646;
or3_6681: n_7637 <=  n_7638  OR n_7641  OR n_7644;
and2_6682: n_7638 <=  n_7639  AND n_7640;
inv_6683: n_7639  <= TRANSPORT NOT a_N2527  ;
delay_6684: n_7640  <= TRANSPORT a_LC6_D5  ;
and2_6685: n_7641 <=  n_7642  AND n_7643;
delay_6686: n_7642  <= TRANSPORT a_N2527  ;
delay_6687: n_7643  <= TRANSPORT a_SCH2BAROUT_F15_G  ;
and1_6688: n_7644 <=  n_7645;
delay_6689: n_7645  <= TRANSPORT a_N818  ;
and1_6690: n_7646 <=  gnd;
delay_6691: n_7647  <= TRANSPORT clk  ;
filter_6692: FILTER_a8237

    PORT MAP (IN1 => n_7647, Y => a_SCH2ADDRREG_F15_G_aCLK);
delay_6693: a_N2555  <= TRANSPORT a_EQ611  ;
xor2_6694: a_EQ611 <=  n_7651  XOR n_7658;
or2_6695: n_7651 <=  n_7652  OR n_7655;
and2_6696: n_7652 <=  n_7653  AND n_7654;
delay_6697: n_7653  <= TRANSPORT a_N2530_aNOT  ;
delay_6698: n_7654  <= TRANSPORT a_N3045  ;
and2_6699: n_7655 <=  n_7656  AND n_7657;
inv_6700: n_7656  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_6701: n_7657  <= TRANSPORT a_SADDRESSOUT_F15_G  ;
and1_6702: n_7658 <=  gnd;
delay_6703: a_LC2_D10  <= TRANSPORT a_EQ649  ;
xor2_6704: a_EQ649 <=  n_7661  XOR n_7673;
or3_6705: n_7661 <=  n_7662  OR n_7666  OR n_7670;
and3_6706: n_7662 <=  n_7663  AND n_7664  AND n_7665;
inv_6707: n_7663  <= TRANSPORT NOT a_LC3_D22  ;
delay_6708: n_7664  <= TRANSPORT a_N2354_aNOT  ;
delay_6709: n_7665  <= TRANSPORT dbin(7)  ;
and2_6710: n_7666 <=  n_7667  AND n_7668;
inv_6711: n_7667  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_6712: n_7668  <= TRANSPORT a_SCH0ADDRREG_F15_G  ;
and2_6713: n_7670 <=  n_7671  AND n_7672;
delay_6714: n_7671  <= TRANSPORT a_LC3_D22  ;
delay_6715: n_7672  <= TRANSPORT a_SCH0ADDRREG_F15_G  ;
and1_6716: n_7673 <=  gnd;
delay_6717: a_LC1_D10  <= TRANSPORT a_EQ650  ;
xor2_6718: a_EQ650 <=  n_7676  XOR n_7683;
or2_6719: n_7676 <=  n_7677  OR n_7680;
and2_6720: n_7677 <=  n_7678  AND n_7679;
inv_6721: n_7678  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_6722: n_7679  <= TRANSPORT a_N2555  ;
and2_6723: n_7680 <=  n_7681  AND n_7682;
delay_6724: n_7681  <= TRANSPORT a_N2558_aNOT  ;
delay_6725: n_7682  <= TRANSPORT a_LC2_D10  ;
and1_6726: n_7683 <=  gnd;
dff_6727: DFF_a8237

    PORT MAP ( D => a_EQ882, CLK => a_SCH0ADDRREG_F15_G_aCLK, CLRN => a_SCH0ADDRREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F15_G);
inv_6728: a_SCH0ADDRREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6729: a_EQ882 <=  n_7690  XOR n_7697;
or2_6730: n_7690 <=  n_7691  OR n_7694;
and2_6731: n_7691 <=  n_7692  AND n_7693;
inv_6732: n_7692  <= TRANSPORT NOT a_N2525  ;
delay_6733: n_7693  <= TRANSPORT a_LC1_D10  ;
and2_6734: n_7694 <=  n_7695  AND n_7696;
delay_6735: n_7695  <= TRANSPORT a_N2525  ;
delay_6736: n_7696  <= TRANSPORT a_SCH0BAROUT_F15_G  ;
and1_6737: n_7697 <=  gnd;
delay_6738: n_7698  <= TRANSPORT clk  ;
filter_6739: FILTER_a8237

    PORT MAP (IN1 => n_7698, Y => a_SCH0ADDRREG_F15_G_aCLK);
delay_6740: a_LC6_D3  <= TRANSPORT a_EQ724  ;
xor2_6741: a_EQ724 <=  n_7702  XOR n_7714;
or3_6742: n_7702 <=  n_7703  OR n_7707  OR n_7711;
and3_6743: n_7703 <=  n_7704  AND n_7705  AND n_7706;
inv_6744: n_7704  <= TRANSPORT NOT a_LC3_D22  ;
inv_6745: n_7705  <= TRANSPORT NOT a_N2348  ;
delay_6746: n_7706  <= TRANSPORT dbin(7)  ;
and2_6747: n_7707 <=  n_7708  AND n_7709;
delay_6748: n_7708  <= TRANSPORT a_N2348  ;
delay_6749: n_7709  <= TRANSPORT a_SCH3ADDRREG_F15_G  ;
and2_6750: n_7711 <=  n_7712  AND n_7713;
delay_6751: n_7712  <= TRANSPORT a_LC3_D22  ;
delay_6752: n_7713  <= TRANSPORT a_SCH3ADDRREG_F15_G  ;
and1_6753: n_7714 <=  gnd;
delay_6754: a_LC5_D3  <= TRANSPORT a_EQ725  ;
xor2_6755: a_EQ725 <=  n_7717  XOR n_7724;
or2_6756: n_7717 <=  n_7718  OR n_7721;
and2_6757: n_7718 <=  n_7719  AND n_7720;
inv_6758: n_7719  <= TRANSPORT NOT a_N965  ;
delay_6759: n_7720  <= TRANSPORT a_N3045  ;
and2_6760: n_7721 <=  n_7722  AND n_7723;
delay_6761: n_7722  <= TRANSPORT a_N965  ;
delay_6762: n_7723  <= TRANSPORT a_LC6_D3  ;
and1_6763: n_7724 <=  gnd;
dff_6764: DFF_a8237

    PORT MAP ( D => a_EQ1074, CLK => a_SCH3ADDRREG_F15_G_aCLK, CLRN => a_SCH3ADDRREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F15_G);
inv_6765: a_SCH3ADDRREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6766: a_EQ1074 <=  n_7731  XOR n_7738;
or2_6767: n_7731 <=  n_7732  OR n_7735;
and2_6768: n_7732 <=  n_7733  AND n_7734;
inv_6769: n_7733  <= TRANSPORT NOT a_N2528  ;
delay_6770: n_7734  <= TRANSPORT a_LC5_D3  ;
and2_6771: n_7735 <=  n_7736  AND n_7737;
delay_6772: n_7736  <= TRANSPORT a_N2528  ;
delay_6773: n_7737  <= TRANSPORT a_SCH3BAROUT_F15_G  ;
and1_6774: n_7738 <=  gnd;
delay_6775: n_7739  <= TRANSPORT clk  ;
filter_6776: FILTER_a8237

    PORT MAP (IN1 => n_7739, Y => a_SCH3ADDRREG_F15_G_aCLK);
delay_6777: a_LC5_D11  <= TRANSPORT a_EQ675  ;
xor2_6778: a_EQ675 <=  n_7743  XOR n_7752;
or2_6779: n_7743 <=  n_7744  OR n_7747;
and2_6780: n_7744 <=  n_7745  AND n_7746;
inv_6781: n_7745  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_6782: n_7746  <= TRANSPORT a_N2555  ;
and3_6783: n_7747 <=  n_7748  AND n_7749  AND n_7750;
delay_6784: n_7748  <= TRANSPORT a_N2585_aNOT  ;
delay_6785: n_7749  <= TRANSPORT a_N2559_aNOT  ;
delay_6786: n_7750  <= TRANSPORT a_SCH1ADDRREG_F15_G  ;
and1_6787: n_7752 <=  gnd;
delay_6788: a_N457  <= TRANSPORT a_N457_aIN  ;
xor2_6789: a_N457_aIN <=  n_7755  XOR n_7761;
or1_6790: n_7755 <=  n_7756;
and4_6791: n_7756 <=  n_7757  AND n_7758  AND n_7759  AND n_7760;
inv_6792: n_7757  <= TRANSPORT NOT a_N2585_aNOT  ;
delay_6793: n_7758  <= TRANSPORT a_N2559_aNOT  ;
inv_6794: n_7759  <= TRANSPORT NOT a_N2526  ;
delay_6795: n_7760  <= TRANSPORT dbin(7)  ;
and1_6796: n_7761 <=  gnd;
dff_6797: DFF_a8237

    PORT MAP ( D => a_EQ946, CLK => a_SCH1ADDRREG_F15_G_aCLK, CLRN => a_SCH1ADDRREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F15_G);
inv_6798: a_SCH1ADDRREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6799: a_EQ946 <=  n_7768  XOR n_7777;
or3_6800: n_7768 <=  n_7769  OR n_7772  OR n_7775;
and2_6801: n_7769 <=  n_7770  AND n_7771;
inv_6802: n_7770  <= TRANSPORT NOT a_N2526  ;
delay_6803: n_7771  <= TRANSPORT a_LC5_D11  ;
and2_6804: n_7772 <=  n_7773  AND n_7774;
delay_6805: n_7773  <= TRANSPORT a_N2526  ;
delay_6806: n_7774  <= TRANSPORT a_SCH1BAROUT_F15_G  ;
and1_6807: n_7775 <=  n_7776;
delay_6808: n_7776  <= TRANSPORT a_N457  ;
and1_6809: n_7777 <=  gnd;
delay_6810: n_7778  <= TRANSPORT clk  ;
filter_6811: FILTER_a8237

    PORT MAP (IN1 => n_7778, Y => a_SCH1ADDRREG_F15_G_aCLK);
delay_6812: a_N63_aNOT  <= TRANSPORT a_EQ184  ;
xor2_6813: a_EQ184 <=  n_7782  XOR n_7791;
or4_6814: n_7782 <=  n_7783  OR n_7785  OR n_7787  OR n_7789;
and1_6815: n_7783 <=  n_7784;
delay_6816: n_7784  <= TRANSPORT ain(2)  ;
and1_6817: n_7785 <=  n_7786;
delay_6818: n_7786  <= TRANSPORT ain(1)  ;
and1_6819: n_7787 <=  n_7788;
inv_6820: n_7788  <= TRANSPORT NOT ain(0)  ;
and1_6821: n_7789 <=  n_7790;
inv_6822: n_7790  <= TRANSPORT NOT ain(3)  ;
and1_6823: n_7791 <=  gnd;
delay_6824: a_N2566_aNOT  <= TRANSPORT a_EQ619  ;
xor2_6825: a_EQ619 <=  n_7794  XOR n_7799;
or2_6826: n_7794 <=  n_7795  OR n_7797;
and1_6827: n_7795 <=  n_7796;
delay_6828: n_7796  <= TRANSPORT a_N63_aNOT  ;
and1_6829: n_7797 <=  n_7798;
delay_6830: n_7798  <= TRANSPORT a_N87  ;
and1_6831: n_7799 <=  gnd;
delay_6832: a_N1434_aNOT  <= TRANSPORT a_EQ439  ;
xor2_6833: a_EQ439 <=  n_7802  XOR n_7812;
or2_6834: n_7802 <=  n_7803  OR n_7808;
and3_6835: n_7803 <=  n_7804  AND n_7805  AND n_7806;
delay_6836: n_7804  <= TRANSPORT a_N2563_aNOT  ;
delay_6837: n_7805  <= TRANSPORT a_N2566_aNOT  ;
delay_6838: n_7806  <= TRANSPORT a_SREQUESTREG_F1_G  ;
and3_6839: n_7808 <=  n_7809  AND n_7810  AND n_7811;
delay_6840: n_7809  <= TRANSPORT a_N2563_aNOT  ;
inv_6841: n_7810  <= TRANSPORT NOT a_N84  ;
delay_6842: n_7811  <= TRANSPORT a_SREQUESTREG_F1_G  ;
and1_6843: n_7812 <=  gnd;
dff_6844: DFF_a8237

    PORT MAP ( D => a_EQ1174, CLK => a_SREQUESTREG_F1_G_aCLK, CLRN => a_SREQUESTREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SREQUESTREG_F1_G);
inv_6845: a_SREQUESTREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6846: a_EQ1174 <=  n_7819  XOR n_7826;
or2_6847: n_7819 <=  n_7820  OR n_7822;
and1_6848: n_7820 <=  n_7821;
delay_6849: n_7821  <= TRANSPORT a_N1434_aNOT  ;
and3_6850: n_7822 <=  n_7823  AND n_7824  AND n_7825;
delay_6851: n_7823  <= TRANSPORT a_N84  ;
inv_6852: n_7824  <= TRANSPORT NOT a_N2566_aNOT  ;
delay_6853: n_7825  <= TRANSPORT dbin(2)  ;
and1_6854: n_7826 <=  gnd;
delay_6855: n_7827  <= TRANSPORT clk  ;
filter_6856: FILTER_a8237

    PORT MAP (IN1 => n_7827, Y => a_SREQUESTREG_F1_G_aCLK);
delay_6857: a_N2582_aNOT  <= TRANSPORT a_EQ634  ;
xor2_6858: a_EQ634 <=  n_7831  XOR n_7836;
or2_6859: n_7831 <=  n_7832  OR n_7834;
and1_6860: n_7832 <=  n_7833;
delay_6861: n_7833  <= TRANSPORT a_N77_aNOT  ;
and1_6862: n_7834 <=  n_7835;
delay_6863: n_7835  <= TRANSPORT a_LC6_D6  ;
and1_6864: n_7836 <=  gnd;
dff_6865: DFF_a8237

    PORT MAP ( D => a_EQ1012, CLK => a_SCH2BAROUT_F1_G_aCLK, CLRN => a_SCH2BAROUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F1_G);
inv_6866: a_SCH2BAROUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6867: a_EQ1012 <=  n_7844  XOR n_7851;
or2_6868: n_7844 <=  n_7845  OR n_7848;
and2_6869: n_7845 <=  n_7846  AND n_7847;
inv_6870: n_7846  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_6871: n_7847  <= TRANSPORT dbin(1)  ;
and2_6872: n_7848 <=  n_7849  AND n_7850;
delay_6873: n_7849  <= TRANSPORT a_N2582_aNOT  ;
delay_6874: n_7850  <= TRANSPORT a_SCH2BAROUT_F1_G  ;
and1_6875: n_7851 <=  gnd;
delay_6876: n_7852  <= TRANSPORT clk  ;
filter_6877: FILTER_a8237

    PORT MAP (IN1 => n_7852, Y => a_SCH2BAROUT_F1_G_aCLK);
delay_6878: a_N2580_aNOT  <= TRANSPORT a_EQ631  ;
xor2_6879: a_EQ631 <=  n_7856  XOR n_7861;
or2_6880: n_7856 <=  n_7857  OR n_7859;
and1_6881: n_7857 <=  n_7858;
delay_6882: n_7858  <= TRANSPORT a_N2348  ;
and1_6883: n_7859 <=  n_7860;
delay_6884: n_7860  <= TRANSPORT a_LC6_D6  ;
and1_6885: n_7861 <=  gnd;
dff_6886: DFF_a8237

    PORT MAP ( D => a_EQ1080, CLK => a_SCH3BAROUT_F5_G_aCLK, CLRN => a_SCH3BAROUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F5_G);
inv_6887: a_SCH3BAROUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6888: a_EQ1080 <=  n_7869  XOR n_7876;
or2_6889: n_7869 <=  n_7870  OR n_7873;
and2_6890: n_7870 <=  n_7871  AND n_7872;
inv_6891: n_7871  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_6892: n_7872  <= TRANSPORT dbin(5)  ;
and2_6893: n_7873 <=  n_7874  AND n_7875;
delay_6894: n_7874  <= TRANSPORT a_N2580_aNOT  ;
delay_6895: n_7875  <= TRANSPORT a_SCH3BAROUT_F5_G  ;
and1_6896: n_7876 <=  gnd;
delay_6897: n_7877  <= TRANSPORT clk  ;
filter_6898: FILTER_a8237

    PORT MAP (IN1 => n_7877, Y => a_SCH3BAROUT_F5_G_aCLK);
dff_6899: DFF_a8237

    PORT MAP ( D => a_EQ1082, CLK => a_SCH3BAROUT_F7_G_aCLK, CLRN => a_SCH3BAROUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F7_G);
inv_6900: a_SCH3BAROUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6901: a_EQ1082 <=  n_7886  XOR n_7893;
or2_6902: n_7886 <=  n_7887  OR n_7890;
and2_6903: n_7887 <=  n_7888  AND n_7889;
inv_6904: n_7888  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_6905: n_7889  <= TRANSPORT dbin(7)  ;
and2_6906: n_7890 <=  n_7891  AND n_7892;
delay_6907: n_7891  <= TRANSPORT a_N2580_aNOT  ;
delay_6908: n_7892  <= TRANSPORT a_SCH3BAROUT_F7_G  ;
and1_6909: n_7893 <=  gnd;
delay_6910: n_7894  <= TRANSPORT clk  ;
filter_6911: FILTER_a8237

    PORT MAP (IN1 => n_7894, Y => a_SCH3BAROUT_F7_G_aCLK);
delay_6912: a_LC3_D21  <= TRANSPORT a_EQ748  ;
xor2_6913: a_EQ748 <=  n_7898  XOR n_7910;
or3_6914: n_7898 <=  n_7899  OR n_7903  OR n_7907;
and3_6915: n_7899 <=  n_7900  AND n_7901  AND n_7902;
inv_6916: n_7900  <= TRANSPORT NOT a_LC3_D22  ;
inv_6917: n_7901  <= TRANSPORT NOT a_N2353  ;
delay_6918: n_7902  <= TRANSPORT dbin(7)  ;
and2_6919: n_7903 <=  n_7904  AND n_7905;
delay_6920: n_7904  <= TRANSPORT a_N2353  ;
delay_6921: n_7905  <= TRANSPORT a_SH0WRDCNTREG_F15_G  ;
and2_6922: n_7907 <=  n_7908  AND n_7909;
delay_6923: n_7908  <= TRANSPORT a_LC3_D22  ;
delay_6924: n_7909  <= TRANSPORT a_SH0WRDCNTREG_F15_G  ;
and1_6925: n_7910 <=  gnd;
delay_6926: a_LC5_D21  <= TRANSPORT a_EQ749  ;
xor2_6927: a_EQ749 <=  n_7913  XOR n_7925;
or3_6928: n_7913 <=  n_7914  OR n_7917  OR n_7921;
and2_6929: n_7914 <=  n_7915  AND n_7916;
delay_6930: n_7915  <= TRANSPORT a_N2558_aNOT  ;
delay_6931: n_7916  <= TRANSPORT a_LC3_D21  ;
and3_6932: n_7917 <=  n_7918  AND n_7919  AND n_7920;
inv_6933: n_7918  <= TRANSPORT NOT a_LC3_E16_aNOT  ;
inv_6934: n_7919  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_6935: n_7920  <= TRANSPORT a_N3541  ;
and3_6936: n_7921 <=  n_7922  AND n_7923  AND n_7924;
delay_6937: n_7922  <= TRANSPORT a_LC3_E16_aNOT  ;
inv_6938: n_7923  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_6939: n_7924  <= TRANSPORT NOT a_N3541  ;
and1_6940: n_7925 <=  gnd;
dff_6941: DFF_a8237

    PORT MAP ( D => a_EQ1138, CLK => a_SH0WRDCNTREG_F15_G_aCLK, CLRN => a_SH0WRDCNTREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SH0WRDCNTREG_F15_G);
inv_6942: a_SH0WRDCNTREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6943: a_EQ1138 <=  n_7932  XOR n_7939;
or2_6944: n_7932 <=  n_7933  OR n_7936;
and2_6945: n_7933 <=  n_7934  AND n_7935;
inv_6946: n_7934  <= TRANSPORT NOT a_N2525  ;
delay_6947: n_7935  <= TRANSPORT a_LC5_D21  ;
and2_6948: n_7936 <=  n_7937  AND n_7938;
delay_6949: n_7937  <= TRANSPORT a_N2525  ;
delay_6950: n_7938  <= TRANSPORT a_SCH0BWORDOUT_F15_G  ;
and1_6951: n_7939 <=  gnd;
delay_6952: n_7940  <= TRANSPORT clk  ;
filter_6953: FILTER_a8237

    PORT MAP (IN1 => n_7940, Y => a_SH0WRDCNTREG_F15_G_aCLK);
delay_6954: a_LC7_D4  <= TRANSPORT a_EQ315  ;
xor2_6955: a_EQ315 <=  n_7944  XOR n_7952;
or2_6956: n_7944 <=  n_7945  OR n_7948;
and2_6957: n_7945 <=  n_7946  AND n_7947;
inv_6958: n_7946  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_6959: n_7947  <= TRANSPORT dbin(7)  ;
and2_6960: n_7948 <=  n_7949  AND n_7950;
delay_6961: n_7949  <= TRANSPORT a_N2577_aNOT  ;
delay_6962: n_7950  <= TRANSPORT a_SH1WRDCNTREG_F15_G  ;
and1_6963: n_7952 <=  gnd;
delay_6964: a_LC5_D4  <= TRANSPORT a_EQ324  ;
xor2_6965: a_EQ324 <=  n_7955  XOR n_7967;
or3_6966: n_7955 <=  n_7956  OR n_7959  OR n_7963;
and2_6967: n_7956 <=  n_7957  AND n_7958;
delay_6968: n_7957  <= TRANSPORT a_N2559_aNOT  ;
delay_6969: n_7958  <= TRANSPORT a_LC7_D4  ;
and3_6970: n_7959 <=  n_7960  AND n_7961  AND n_7962;
inv_6971: n_7960  <= TRANSPORT NOT a_LC3_E16_aNOT  ;
inv_6972: n_7961  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_6973: n_7962  <= TRANSPORT a_N3541  ;
and3_6974: n_7963 <=  n_7964  AND n_7965  AND n_7966;
delay_6975: n_7964  <= TRANSPORT a_LC3_E16_aNOT  ;
inv_6976: n_7965  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_6977: n_7966  <= TRANSPORT NOT a_N3541  ;
and1_6978: n_7967 <=  gnd;
dff_6979: DFF_a8237

    PORT MAP ( D => a_EQ1144, CLK => a_SH1WRDCNTREG_F15_G_aCLK, CLRN => a_SH1WRDCNTREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SH1WRDCNTREG_F15_G);
inv_6980: a_SH1WRDCNTREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_6981: a_EQ1144 <=  n_7974  XOR n_7981;
or2_6982: n_7974 <=  n_7975  OR n_7978;
and2_6983: n_7975 <=  n_7976  AND n_7977;
inv_6984: n_7976  <= TRANSPORT NOT a_N2526  ;
delay_6985: n_7977  <= TRANSPORT a_LC5_D4  ;
and2_6986: n_7978 <=  n_7979  AND n_7980;
delay_6987: n_7979  <= TRANSPORT a_N2526  ;
delay_6988: n_7980  <= TRANSPORT a_SCH1BWORDOUT_F15_G  ;
and1_6989: n_7981 <=  gnd;
delay_6990: n_7982  <= TRANSPORT clk  ;
filter_6991: FILTER_a8237

    PORT MAP (IN1 => n_7982, Y => a_SH1WRDCNTREG_F15_G_aCLK);
delay_6992: a_N1149_aNOT  <= TRANSPORT a_EQ370  ;
xor2_6993: a_EQ370 <=  n_7986  XOR n_7998;
or3_6994: n_7986 <=  n_7987  OR n_7991  OR n_7995;
and3_6995: n_7987 <=  n_7988  AND n_7989  AND n_7990;
inv_6996: n_7988  <= TRANSPORT NOT a_LC3_D22  ;
inv_6997: n_7989  <= TRANSPORT NOT a_N62_aNOT  ;
delay_6998: n_7990  <= TRANSPORT dbin(7)  ;
and2_6999: n_7991 <=  n_7992  AND n_7993;
delay_7000: n_7992  <= TRANSPORT a_N62_aNOT  ;
delay_7001: n_7993  <= TRANSPORT a_SH2WRDCNTREG_F15_G  ;
and2_7002: n_7995 <=  n_7996  AND n_7997;
delay_7003: n_7996  <= TRANSPORT a_LC3_D22  ;
delay_7004: n_7997  <= TRANSPORT a_SH2WRDCNTREG_F15_G  ;
and1_7005: n_7998 <=  gnd;
delay_7006: a_LC1_D7  <= TRANSPORT a_EQ371  ;
xor2_7007: a_EQ371 <=  n_8001  XOR n_8013;
or3_7008: n_8001 <=  n_8002  OR n_8005  OR n_8009;
and2_7009: n_8002 <=  n_8003  AND n_8004;
delay_7010: n_8003  <= TRANSPORT a_N2560_aNOT  ;
delay_7011: n_8004  <= TRANSPORT a_N1149_aNOT  ;
and3_7012: n_8005 <=  n_8006  AND n_8007  AND n_8008;
inv_7013: n_8006  <= TRANSPORT NOT a_LC3_E16_aNOT  ;
inv_7014: n_8007  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_7015: n_8008  <= TRANSPORT a_N3541  ;
and3_7016: n_8009 <=  n_8010  AND n_8011  AND n_8012;
delay_7017: n_8010  <= TRANSPORT a_LC3_E16_aNOT  ;
inv_7018: n_8011  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_7019: n_8012  <= TRANSPORT NOT a_N3541  ;
and1_7020: n_8013 <=  gnd;
dff_7021: DFF_a8237

    PORT MAP ( D => a_EQ1150, CLK => a_SH2WRDCNTREG_F15_G_aCLK, CLRN => a_SH2WRDCNTREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SH2WRDCNTREG_F15_G);
inv_7022: a_SH2WRDCNTREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7023: a_EQ1150 <=  n_8020  XOR n_8027;
or2_7024: n_8020 <=  n_8021  OR n_8024;
and2_7025: n_8021 <=  n_8022  AND n_8023;
delay_7026: n_8022  <= TRANSPORT a_N2527  ;
delay_7027: n_8023  <= TRANSPORT a_SCH2BWORDOUT_F15_G  ;
and2_7028: n_8024 <=  n_8025  AND n_8026;
inv_7029: n_8025  <= TRANSPORT NOT a_N2527  ;
delay_7030: n_8026  <= TRANSPORT a_LC1_D7  ;
and1_7031: n_8027 <=  gnd;
delay_7032: n_8028  <= TRANSPORT clk  ;
filter_7033: FILTER_a8237

    PORT MAP (IN1 => n_8028, Y => a_SH2WRDCNTREG_F15_G_aCLK);
delay_7034: a_LC2_D3  <= TRANSPORT a_EQ814  ;
xor2_7035: a_EQ814 <=  n_8032  XOR n_8040;
or2_7036: n_8032 <=  n_8033  OR n_8036;
and2_7037: n_8033 <=  n_8034  AND n_8035;
inv_7038: n_8034  <= TRANSPORT NOT a_N2573_aNOT  ;
delay_7039: n_8035  <= TRANSPORT dbin(7)  ;
and2_7040: n_8036 <=  n_8037  AND n_8038;
delay_7041: n_8037  <= TRANSPORT a_N2573_aNOT  ;
delay_7042: n_8038  <= TRANSPORT a_SH3WRDCNTREG_F15_G  ;
and1_7043: n_8040 <=  gnd;
delay_7044: a_LC3_D3  <= TRANSPORT a_EQ815  ;
xor2_7045: a_EQ815 <=  n_8043  XOR n_8055;
or3_7046: n_8043 <=  n_8044  OR n_8047  OR n_8051;
and2_7047: n_8044 <=  n_8045  AND n_8046;
delay_7048: n_8045  <= TRANSPORT a_N965  ;
delay_7049: n_8046  <= TRANSPORT a_LC2_D3  ;
and3_7050: n_8047 <=  n_8048  AND n_8049  AND n_8050;
inv_7051: n_8048  <= TRANSPORT NOT a_LC3_E16_aNOT  ;
inv_7052: n_8049  <= TRANSPORT NOT a_N965  ;
delay_7053: n_8050  <= TRANSPORT a_N3541  ;
and3_7054: n_8051 <=  n_8052  AND n_8053  AND n_8054;
delay_7055: n_8052  <= TRANSPORT a_LC3_E16_aNOT  ;
inv_7056: n_8053  <= TRANSPORT NOT a_N965  ;
inv_7057: n_8054  <= TRANSPORT NOT a_N3541  ;
and1_7058: n_8055 <=  gnd;
dff_7059: DFF_a8237

    PORT MAP ( D => a_EQ1156, CLK => a_SH3WRDCNTREG_F15_G_aCLK, CLRN => a_SH3WRDCNTREG_F15_G_aCLRN,
          PRN => vcc, Q => a_SH3WRDCNTREG_F15_G);
inv_7060: a_SH3WRDCNTREG_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7061: a_EQ1156 <=  n_8062  XOR n_8069;
or2_7062: n_8062 <=  n_8063  OR n_8066;
and2_7063: n_8063 <=  n_8064  AND n_8065;
inv_7064: n_8064  <= TRANSPORT NOT a_N2528  ;
delay_7065: n_8065  <= TRANSPORT a_LC3_D3  ;
and2_7066: n_8066 <=  n_8067  AND n_8068;
delay_7067: n_8067  <= TRANSPORT a_N2528  ;
delay_7068: n_8068  <= TRANSPORT a_SCH3BWORDOUT_F15_G  ;
and1_7069: n_8069 <=  gnd;
delay_7070: n_8070  <= TRANSPORT clk  ;
filter_7071: FILTER_a8237

    PORT MAP (IN1 => n_8070, Y => a_SH3WRDCNTREG_F15_G_aCLK);
delay_7072: a_LC2_D24  <= TRANSPORT a_EQ277  ;
xor2_7073: a_EQ277 <=  n_8074  XOR n_8085;
or3_7074: n_8074 <=  n_8075  OR n_8078  OR n_8081;
and2_7075: n_8075 <=  n_8076  AND n_8077;
inv_7076: n_8076  <= TRANSPORT NOT a_LC8_F13_aNOT  ;
delay_7077: n_8077  <= TRANSPORT a_N3549  ;
and2_7078: n_8078 <=  n_8079  AND n_8080;
inv_7079: n_8079  <= TRANSPORT NOT a_N2557  ;
delay_7080: n_8080  <= TRANSPORT a_N3549  ;
and3_7081: n_8081 <=  n_8082  AND n_8083  AND n_8084;
delay_7082: n_8082  <= TRANSPORT a_N2557  ;
delay_7083: n_8083  <= TRANSPORT a_LC8_F13_aNOT  ;
inv_7084: n_8084  <= TRANSPORT NOT a_N3549  ;
and1_7085: n_8085 <=  gnd;
delay_7086: a_LC4_D24  <= TRANSPORT a_EQ276  ;
xor2_7087: a_EQ276 <=  n_8088  XOR n_8095;
or2_7088: n_8088 <=  n_8089  OR n_8092;
and2_7089: n_8089 <=  n_8090  AND n_8091;
delay_7090: n_8090  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_7091: n_8091  <= TRANSPORT a_SCH1WRDCNTREG_F7_G  ;
and2_7092: n_8092 <=  n_8093  AND n_8094;
inv_7093: n_8093  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_7094: n_8094  <= TRANSPORT a_SCH0WRDCNTREG_F7_G  ;
and1_7095: n_8095 <=  gnd;
delay_7096: a_N629_aNOT  <= TRANSPORT a_EQ274  ;
xor2_7097: a_EQ274 <=  n_8098  XOR n_8105;
or2_7098: n_8098 <=  n_8099  OR n_8102;
and2_7099: n_8099 <=  n_8100  AND n_8101;
inv_7100: n_8100  <= TRANSPORT NOT a_N2531  ;
delay_7101: n_8101  <= TRANSPORT a_LC2_D24  ;
and2_7102: n_8102 <=  n_8103  AND n_8104;
delay_7103: n_8103  <= TRANSPORT a_N2531  ;
delay_7104: n_8104  <= TRANSPORT a_LC4_D24  ;
and1_7105: n_8105 <=  gnd;
delay_7106: a_LC4_D15  <= TRANSPORT a_EQ273  ;
xor2_7107: a_EQ273 <=  n_8108  XOR n_8115;
or2_7108: n_8108 <=  n_8109  OR n_8112;
and2_7109: n_8109 <=  n_8110  AND n_8111;
inv_7110: n_8110  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_7111: n_8111  <= TRANSPORT a_SCH0WRDCNTREG_F7_G  ;
and2_7112: n_8112 <=  n_8113  AND n_8114;
inv_7113: n_8113  <= TRANSPORT NOT a_N88_aNOT  ;
delay_7114: n_8114  <= TRANSPORT a_SCH1WRDCNTREG_F7_G  ;
and1_7115: n_8115 <=  gnd;
delay_7116: a_LC2_D15  <= TRANSPORT a_EQ272  ;
xor2_7117: a_EQ272 <=  n_8118  XOR n_8125;
or2_7118: n_8118 <=  n_8119  OR n_8122;
and2_7119: n_8119 <=  n_8120  AND n_8121;
inv_7120: n_8120  <= TRANSPORT NOT a_N2377  ;
delay_7121: n_8121  <= TRANSPORT a_SCH3WRDCNTREG_F7_G  ;
and2_7122: n_8122 <=  n_8123  AND n_8124;
inv_7123: n_8123  <= TRANSPORT NOT a_N2376  ;
delay_7124: n_8124  <= TRANSPORT a_SCH2WRDCNTREG_F7_G  ;
and1_7125: n_8125 <=  gnd;
dff_7126: DFF_a8237

    PORT MAP ( D => a_EQ845, CLK => a_N3549_aCLK, CLRN => a_N3549_aCLRN, PRN => vcc,
          Q => a_N3549);
inv_7127: a_N3549_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7128: a_EQ845 <=  n_8132  XOR n_8142;
or3_7129: n_8132 <=  n_8133  OR n_8136  OR n_8139;
and2_7130: n_8133 <=  n_8134  AND n_8135;
delay_7131: n_8134  <= TRANSPORT a_N629_aNOT  ;
inv_7132: n_8135  <= TRANSPORT NOT startdma  ;
and2_7133: n_8136 <=  n_8137  AND n_8138;
delay_7134: n_8137  <= TRANSPORT a_LC4_D15  ;
delay_7135: n_8138  <= TRANSPORT startdma  ;
and2_7136: n_8139 <=  n_8140  AND n_8141;
delay_7137: n_8140  <= TRANSPORT a_LC2_D15  ;
delay_7138: n_8141  <= TRANSPORT startdma  ;
and1_7139: n_8142 <=  gnd;
delay_7140: n_8143  <= TRANSPORT clk  ;
filter_7141: FILTER_a8237

    PORT MAP (IN1 => n_8143, Y => a_N3549_aCLK);
delay_7142: a_N1174  <= TRANSPORT a_EQ381  ;
xor2_7143: a_EQ381 <=  n_8147  XOR n_8154;
or2_7144: n_8147 <=  n_8148  OR n_8151;
and2_7145: n_8148 <=  n_8149  AND n_8150;
inv_7146: n_8149  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_7147: n_8150  <= TRANSPORT a_SCH0WRDCNTREG_F8_G  ;
and2_7148: n_8151 <=  n_8152  AND n_8153;
delay_7149: n_8152  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_7150: n_8153  <= TRANSPORT a_SCH1WRDCNTREG_F8_G  ;
and1_7151: n_8154 <=  gnd;
delay_7152: a_N1163_aNOT  <= TRANSPORT a_EQ373  ;
xor2_7153: a_EQ373 <=  n_8157  XOR n_8164;
or2_7154: n_8157 <=  n_8158  OR n_8161;
and2_7155: n_8158 <=  n_8159  AND n_8160;
inv_7156: n_8159  <= TRANSPORT NOT a_N2557  ;
delay_7157: n_8160  <= TRANSPORT a_N3548  ;
and2_7158: n_8161 <=  n_8162  AND n_8163;
delay_7159: n_8162  <= TRANSPORT a_N2557  ;
inv_7160: n_8163  <= TRANSPORT NOT a_LC6_D17  ;
and1_7161: n_8164 <=  gnd;
delay_7162: a_LC6_D24  <= TRANSPORT a_EQ382  ;
xor2_7163: a_EQ382 <=  n_8167  XOR n_8174;
or2_7164: n_8167 <=  n_8168  OR n_8171;
and2_7165: n_8168 <=  n_8169  AND n_8170;
delay_7166: n_8169  <= TRANSPORT a_N2531  ;
delay_7167: n_8170  <= TRANSPORT a_N1174  ;
and2_7168: n_8171 <=  n_8172  AND n_8173;
inv_7169: n_8172  <= TRANSPORT NOT a_N2531  ;
delay_7170: n_8173  <= TRANSPORT a_N1163_aNOT  ;
and1_7171: n_8174 <=  gnd;
delay_7172: a_LC1_D6  <= TRANSPORT a_EQ380  ;
xor2_7173: a_EQ380 <=  n_8177  XOR n_8184;
or2_7174: n_8177 <=  n_8178  OR n_8181;
and2_7175: n_8178 <=  n_8179  AND n_8180;
inv_7176: n_8179  <= TRANSPORT NOT a_N88_aNOT  ;
delay_7177: n_8180  <= TRANSPORT a_SCH1WRDCNTREG_F8_G  ;
and2_7178: n_8181 <=  n_8182  AND n_8183;
inv_7179: n_8182  <= TRANSPORT NOT a_N2377  ;
delay_7180: n_8183  <= TRANSPORT a_SCH3WRDCNTREG_F8_G  ;
and1_7181: n_8184 <=  gnd;
delay_7182: a_LC1_D24  <= TRANSPORT a_EQ379  ;
xor2_7183: a_EQ379 <=  n_8187  XOR n_8194;
or2_7184: n_8187 <=  n_8188  OR n_8191;
and2_7185: n_8188 <=  n_8189  AND n_8190;
inv_7186: n_8189  <= TRANSPORT NOT a_N2376  ;
delay_7187: n_8190  <= TRANSPORT a_SCH2WRDCNTREG_F8_G  ;
and2_7188: n_8191 <=  n_8192  AND n_8193;
inv_7189: n_8192  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_7190: n_8193  <= TRANSPORT a_SCH0WRDCNTREG_F8_G  ;
and1_7191: n_8194 <=  gnd;
dff_7192: DFF_a8237

    PORT MAP ( D => a_EQ844, CLK => a_N3548_aCLK, CLRN => a_N3548_aCLRN, PRN => vcc,
          Q => a_N3548);
inv_7193: a_N3548_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7194: a_EQ844 <=  n_8201  XOR n_8211;
or3_7195: n_8201 <=  n_8202  OR n_8205  OR n_8208;
and2_7196: n_8202 <=  n_8203  AND n_8204;
delay_7197: n_8203  <= TRANSPORT a_LC6_D24  ;
inv_7198: n_8204  <= TRANSPORT NOT startdma  ;
and2_7199: n_8205 <=  n_8206  AND n_8207;
delay_7200: n_8206  <= TRANSPORT a_LC1_D6  ;
delay_7201: n_8207  <= TRANSPORT startdma  ;
and2_7202: n_8208 <=  n_8209  AND n_8210;
delay_7203: n_8209  <= TRANSPORT a_LC1_D24  ;
delay_7204: n_8210  <= TRANSPORT startdma  ;
and1_7205: n_8211 <=  gnd;
delay_7206: n_8212  <= TRANSPORT clk  ;
filter_7207: FILTER_a8237

    PORT MAP (IN1 => n_8212, Y => a_N3548_aCLK);
delay_7208: a_LC5_A13  <= TRANSPORT a_EQ227  ;
xor2_7209: a_EQ227 <=  n_8216  XOR n_8223;
or2_7210: n_8216 <=  n_8217  OR n_8220;
and2_7211: n_8217 <=  n_8218  AND n_8219;
delay_7212: n_8218  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_7213: n_8219  <= TRANSPORT a_SCH1WRDCNTREG_F9_G  ;
and2_7214: n_8220 <=  n_8221  AND n_8222;
inv_7215: n_8221  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_7216: n_8222  <= TRANSPORT a_SCH0WRDCNTREG_F9_G  ;
and1_7217: n_8223 <=  gnd;
delay_7218: a_LC2_A13  <= TRANSPORT a_EQ225  ;
xor2_7219: a_EQ225 <=  n_8226  XOR n_8236;
or3_7220: n_8226 <=  n_8227  OR n_8230  OR n_8233;
and2_7221: n_8227 <=  n_8228  AND n_8229;
delay_7222: n_8228  <= TRANSPORT a_N2557  ;
inv_7223: n_8229  <= TRANSPORT NOT a_LC1_A13  ;
and2_7224: n_8230 <=  n_8231  AND n_8232;
delay_7225: n_8231  <= TRANSPORT a_N2557  ;
delay_7226: n_8232  <= TRANSPORT a_N2531  ;
and2_7227: n_8233 <=  n_8234  AND n_8235;
inv_7228: n_8234  <= TRANSPORT NOT a_N2557  ;
delay_7229: n_8235  <= TRANSPORT a_N3547  ;
and1_7230: n_8236 <=  gnd;
delay_7231: a_N295_aNOT  <= TRANSPORT a_EQ226  ;
xor2_7232: a_EQ226 <=  n_8239  XOR n_8246;
or2_7233: n_8239 <=  n_8240  OR n_8243;
and2_7234: n_8240 <=  n_8241  AND n_8242;
delay_7235: n_8241  <= TRANSPORT a_LC5_A13  ;
delay_7236: n_8242  <= TRANSPORT a_LC2_A13  ;
and2_7237: n_8243 <=  n_8244  AND n_8245;
inv_7238: n_8244  <= TRANSPORT NOT a_N2531  ;
delay_7239: n_8245  <= TRANSPORT a_LC2_A13  ;
and1_7240: n_8246 <=  gnd;
delay_7241: a_LC8_A13  <= TRANSPORT a_EQ229  ;
xor2_7242: a_EQ229 <=  n_8249  XOR n_8256;
or2_7243: n_8249 <=  n_8250  OR n_8253;
and2_7244: n_8250 <=  n_8251  AND n_8252;
inv_7245: n_8251  <= TRANSPORT NOT a_N2377  ;
delay_7246: n_8252  <= TRANSPORT a_SCH3WRDCNTREG_F9_G  ;
and2_7247: n_8253 <=  n_8254  AND n_8255;
inv_7248: n_8254  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_7249: n_8255  <= TRANSPORT a_SCH0WRDCNTREG_F9_G  ;
and1_7250: n_8256 <=  gnd;
delay_7251: a_LC7_A13  <= TRANSPORT a_EQ228  ;
xor2_7252: a_EQ228 <=  n_8259  XOR n_8266;
or2_7253: n_8259 <=  n_8260  OR n_8263;
and2_7254: n_8260 <=  n_8261  AND n_8262;
inv_7255: n_8261  <= TRANSPORT NOT a_N2376  ;
delay_7256: n_8262  <= TRANSPORT a_SCH2WRDCNTREG_F9_G  ;
and2_7257: n_8263 <=  n_8264  AND n_8265;
inv_7258: n_8264  <= TRANSPORT NOT a_N88_aNOT  ;
delay_7259: n_8265  <= TRANSPORT a_SCH1WRDCNTREG_F9_G  ;
and1_7260: n_8266 <=  gnd;
dff_7261: DFF_a8237

    PORT MAP ( D => a_EQ843, CLK => a_N3547_aCLK, CLRN => a_N3547_aCLRN, PRN => vcc,
          Q => a_N3547);
inv_7262: a_N3547_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7263: a_EQ843 <=  n_8273  XOR n_8283;
or3_7264: n_8273 <=  n_8274  OR n_8277  OR n_8280;
and2_7265: n_8274 <=  n_8275  AND n_8276;
delay_7266: n_8275  <= TRANSPORT a_N295_aNOT  ;
inv_7267: n_8276  <= TRANSPORT NOT startdma  ;
and2_7268: n_8277 <=  n_8278  AND n_8279;
delay_7269: n_8278  <= TRANSPORT a_LC8_A13  ;
delay_7270: n_8279  <= TRANSPORT startdma  ;
and2_7271: n_8280 <=  n_8281  AND n_8282;
delay_7272: n_8281  <= TRANSPORT a_LC7_A13  ;
delay_7273: n_8282  <= TRANSPORT startdma  ;
and1_7274: n_8283 <=  gnd;
delay_7275: n_8284  <= TRANSPORT clk  ;
filter_7276: FILTER_a8237

    PORT MAP (IN1 => n_8284, Y => a_N3547_aCLK);
delay_7277: a_N73  <= TRANSPORT a_N73_aIN  ;
xor2_7278: a_N73_aIN <=  n_8288  XOR n_8294;
or1_7279: n_8288 <=  n_8289;
and4_7280: n_8289 <=  n_8290  AND n_8291  AND n_8292  AND n_8293;
delay_7281: n_8290  <= TRANSPORT ain(3)  ;
inv_7282: n_8291  <= TRANSPORT NOT ain(2)  ;
delay_7283: n_8292  <= TRANSPORT ain(1)  ;
inv_7284: n_8293  <= TRANSPORT NOT ain(0)  ;
and1_7285: n_8294 <=  gnd;
delay_7286: a_N65  <= TRANSPORT a_N65_aIN  ;
xor2_7287: a_N65_aIN <=  n_8297  XOR n_8303;
or1_7288: n_8297 <=  n_8298;
and4_7289: n_8298 <=  n_8299  AND n_8300  AND n_8301  AND n_8302;
delay_7290: n_8299  <= TRANSPORT ain(3)  ;
delay_7291: n_8300  <= TRANSPORT ain(2)  ;
delay_7292: n_8301  <= TRANSPORT ain(1)  ;
delay_7293: n_8302  <= TRANSPORT ain(0)  ;
and1_7294: n_8303 <=  gnd;
delay_7295: a_N1119_aNOT  <= TRANSPORT a_EQ359  ;
xor2_7296: a_EQ359 <=  n_8306  XOR n_8312;
or2_7297: n_8306 <=  n_8307  OR n_8310;
and2_7298: n_8307 <=  n_8308  AND n_8309;
inv_7299: n_8308  <= TRANSPORT NOT a_N73  ;
inv_7300: n_8309  <= TRANSPORT NOT a_N65  ;
and1_7301: n_8310 <=  n_8311;
delay_7302: n_8311  <= TRANSPORT a_N87  ;
and1_7303: n_8312 <=  gnd;
delay_7304: a_N1103_aNOT  <= TRANSPORT a_EQ354  ;
xor2_7305: a_EQ354 <=  n_8315  XOR n_8325;
or2_7306: n_8315 <=  n_8316  OR n_8321;
and3_7307: n_8316 <=  n_8317  AND n_8318  AND n_8319;
inv_7308: n_8317  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7309: n_8318  <= TRANSPORT a_N1119_aNOT  ;
delay_7310: n_8319  <= TRANSPORT a_SMASKREG_F0_G_aNOT  ;
and3_7311: n_8321 <=  n_8322  AND n_8323  AND n_8324;
delay_7312: n_8322  <= TRANSPORT a_N2598_aNOT  ;
delay_7313: n_8323  <= TRANSPORT a_N1119_aNOT  ;
delay_7314: n_8324  <= TRANSPORT a_SMASKREG_F0_G_aNOT  ;
and1_7315: n_8325 <=  gnd;
delay_7316: a_N2564  <= TRANSPORT a_N2564_aIN  ;
xor2_7317: a_N2564_aIN <=  n_8328  XOR n_8332;
or1_7318: n_8328 <=  n_8329;
and2_7319: n_8329 <=  n_8330  AND n_8331;
inv_7320: n_8330  <= TRANSPORT NOT a_N87  ;
delay_7321: n_8331  <= TRANSPORT a_N65  ;
and1_7322: n_8332 <=  gnd;
delay_7323: a_LC2_B4_aNOT  <= TRANSPORT a_EQ356  ;
xor2_7324: a_EQ356 <=  n_8335  XOR n_8343;
or2_7325: n_8335 <=  n_8336  OR n_8340;
and3_7326: n_8336 <=  n_8337  AND n_8338  AND n_8339;
delay_7327: n_8337  <= TRANSPORT a_N2598_aNOT  ;
delay_7328: n_8338  <= TRANSPORT a_N2564  ;
delay_7329: n_8339  <= TRANSPORT a_SMASKREG_F0_G_aNOT  ;
and2_7330: n_8340 <=  n_8341  AND n_8342;
inv_7331: n_8341  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_7332: n_8342  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and1_7333: n_8343 <=  gnd;
delay_7334: a_N75_aNOT  <= TRANSPORT a_EQ193  ;
xor2_7335: a_EQ193 <=  n_8346  XOR n_8355;
or4_7336: n_8346 <=  n_8347  OR n_8349  OR n_8351  OR n_8353;
and1_7337: n_8347 <=  n_8348;
inv_7338: n_8348  <= TRANSPORT NOT ain(2)  ;
and1_7339: n_8349 <=  n_8350;
inv_7340: n_8350  <= TRANSPORT NOT ain(1)  ;
and1_7341: n_8351 <=  n_8352;
delay_7342: n_8352  <= TRANSPORT ain(0)  ;
and1_7343: n_8353 <=  n_8354;
inv_7344: n_8354  <= TRANSPORT NOT ain(3)  ;
and1_7345: n_8355 <=  gnd;
delay_7346: a_N103_aNOT  <= TRANSPORT a_N103_aNOT_aIN  ;
xor2_7347: a_N103_aNOT_aIN <=  n_8358  XOR n_8362;
or1_7348: n_8358 <=  n_8359;
and2_7349: n_8359 <=  n_8360  AND n_8361;
inv_7350: n_8360  <= TRANSPORT NOT a_N87  ;
inv_7351: n_8361  <= TRANSPORT NOT a_N75_aNOT  ;
and1_7352: n_8362 <=  gnd;
delay_7353: a_LC1_B4  <= TRANSPORT a_EQ357  ;
xor2_7354: a_EQ357 <=  n_8365  XOR n_8371;
or2_7355: n_8365 <=  n_8366  OR n_8369;
and2_7356: n_8366 <=  n_8367  AND n_8368;
delay_7357: n_8367  <= TRANSPORT a_N57_aNOT  ;
delay_7358: n_8368  <= TRANSPORT a_LC2_B4_aNOT  ;
and1_7359: n_8369 <=  n_8370;
delay_7360: n_8370  <= TRANSPORT a_N103_aNOT  ;
and1_7361: n_8371 <=  gnd;
delay_7362: a_N104_aNOT  <= TRANSPORT a_N104_aNOT_aIN  ;
xor2_7363: a_N104_aNOT_aIN <=  n_8374  XOR n_8378;
or1_7364: n_8374 <=  n_8375;
and2_7365: n_8375 <=  n_8376  AND n_8377;
inv_7366: n_8376  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7367: n_8377  <= TRANSPORT a_N2564  ;
and1_7368: n_8378 <=  gnd;
delay_7369: a_LC7_B4  <= TRANSPORT a_EQ358  ;
xor2_7370: a_EQ358 <=  n_8381  XOR n_8389;
or3_7371: n_8381 <=  n_8382  OR n_8384  OR n_8386;
and1_7372: n_8382 <=  n_8383;
delay_7373: n_8383  <= TRANSPORT a_N1103_aNOT  ;
and1_7374: n_8384 <=  n_8385;
delay_7375: n_8385  <= TRANSPORT a_LC1_B4  ;
and2_7376: n_8386 <=  n_8387  AND n_8388;
delay_7377: n_8387  <= TRANSPORT a_N104_aNOT  ;
inv_7378: n_8388  <= TRANSPORT NOT dbin(0)  ;
and1_7379: n_8389 <=  gnd;
delay_7380: a_LC5_B4_aNOT  <= TRANSPORT a_EQ353  ;
xor2_7381: a_EQ353 <=  n_8392  XOR n_8399;
or2_7382: n_8392 <=  n_8393  OR n_8396;
and2_7383: n_8393 <=  n_8394  AND n_8395;
inv_7384: n_8394  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7385: n_8395  <= TRANSPORT a_SMASKREG_F0_G_aNOT  ;
and2_7386: n_8396 <=  n_8397  AND n_8398;
delay_7387: n_8397  <= TRANSPORT a_N2598_aNOT  ;
delay_7388: n_8398  <= TRANSPORT a_SMASKREG_F0_G_aNOT  ;
and1_7389: n_8399 <=  gnd;
delay_7390: a_N1108  <= TRANSPORT a_EQ355  ;
xor2_7391: a_EQ355 <=  n_8402  XOR n_8413;
or3_7392: n_8402 <=  n_8403  OR n_8406  OR n_8409;
and2_7393: n_8403 <=  n_8404  AND n_8405;
inv_7394: n_8404  <= TRANSPORT NOT a_N2532_aNOT  ;
delay_7395: n_8405  <= TRANSPORT a_LC5_B4_aNOT  ;
and2_7396: n_8406 <=  n_8407  AND n_8408;
delay_7397: n_8407  <= TRANSPORT a_N57_aNOT  ;
delay_7398: n_8408  <= TRANSPORT a_LC5_B4_aNOT  ;
and3_7399: n_8409 <=  n_8410  AND n_8411  AND n_8412;
inv_7400: n_8410  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7401: n_8411  <= TRANSPORT a_N2532_aNOT  ;
inv_7402: n_8412  <= TRANSPORT NOT dbin(2)  ;
and1_7403: n_8413 <=  gnd;
delay_7404: a_N2565  <= TRANSPORT a_N2565_aIN  ;
xor2_7405: a_N2565_aIN <=  n_8416  XOR n_8420;
or1_7406: n_8416 <=  n_8417;
and2_7407: n_8417 <=  n_8418  AND n_8419;
inv_7408: n_8418  <= TRANSPORT NOT a_N87  ;
delay_7409: n_8419  <= TRANSPORT a_N73  ;
and1_7410: n_8420 <=  gnd;
dff_7411: DFF_a8237

    PORT MAP ( D => a_EQ1157, CLK => a_SMASKREG_F0_G_aNOT_aCLK, CLRN => a_SMASKREG_F0_G_aNOT_aCLRN,
          PRN => vcc, Q => a_SMASKREG_F0_G_aNOT);
inv_7412: a_SMASKREG_F0_G_aNOT_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7413: a_EQ1157 <=  n_8427  XOR n_8435;
or2_7414: n_8427 <=  n_8428  OR n_8431;
and2_7415: n_8428 <=  n_8429  AND n_8430;
delay_7416: n_8429  <= TRANSPORT a_N2563_aNOT  ;
delay_7417: n_8430  <= TRANSPORT a_LC7_B4  ;
and3_7418: n_8431 <=  n_8432  AND n_8433  AND n_8434;
delay_7419: n_8432  <= TRANSPORT a_N2563_aNOT  ;
delay_7420: n_8433  <= TRANSPORT a_N1108  ;
delay_7421: n_8434  <= TRANSPORT a_N2565  ;
and1_7422: n_8435 <=  gnd;
delay_7423: n_8436  <= TRANSPORT clk  ;
filter_7424: FILTER_a8237

    PORT MAP (IN1 => n_8436, Y => a_SMASKREG_F0_G_aNOT_aCLK);
delay_7425: a_N45  <= TRANSPORT a_N45_aIN  ;
xor2_7426: a_N45_aIN <=  n_8440  XOR n_8445;
or1_7427: n_8440 <=  n_8441;
and3_7428: n_8441 <=  n_8442  AND n_8443  AND n_8444;
inv_7429: n_8442  <= TRANSPORT NOT a_N87  ;
delay_7430: n_8443  <= TRANSPORT a_N2532_aNOT  ;
inv_7431: n_8444  <= TRANSPORT NOT a_N63_aNOT  ;
and1_7432: n_8445 <=  gnd;
dff_7433: DFF_a8237

    PORT MAP ( D => a_EQ1173, CLK => a_SREQUESTREG_F0_G_aCLK, CLRN => a_SREQUESTREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SREQUESTREG_F0_G);
inv_7434: a_SREQUESTREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7435: a_EQ1173 <=  n_8453  XOR n_8462;
or2_7436: n_8453 <=  n_8454  OR n_8458;
and3_7437: n_8454 <=  n_8455  AND n_8456  AND n_8457;
delay_7438: n_8455  <= TRANSPORT a_N2563_aNOT  ;
inv_7439: n_8456  <= TRANSPORT NOT a_N45  ;
delay_7440: n_8457  <= TRANSPORT a_SREQUESTREG_F0_G  ;
and3_7441: n_8458 <=  n_8459  AND n_8460  AND n_8461;
delay_7442: n_8459  <= TRANSPORT a_N2563_aNOT  ;
delay_7443: n_8460  <= TRANSPORT a_N45  ;
delay_7444: n_8461  <= TRANSPORT dbin(2)  ;
and1_7445: n_8462 <=  gnd;
delay_7446: n_8463  <= TRANSPORT clk  ;
filter_7447: FILTER_a8237

    PORT MAP (IN1 => n_8463, Y => a_SREQUESTREG_F0_G_aCLK);
delay_7448: a_N1530_aNOT  <= TRANSPORT a_EQ458  ;
xor2_7449: a_EQ458 <=  n_8467  XOR n_8475;
or2_7450: n_8467 <=  n_8468  OR n_8471;
and1_7451: n_8468 <=  n_8469;
delay_7452: n_8469  <= TRANSPORT a_STCSTATUS_F0_G  ;
and3_7453: n_8471 <=  n_8472  AND n_8473  AND n_8474;
inv_7454: n_8472  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_7455: n_8473  <= TRANSPORT a_N57_aNOT  ;
inv_7456: n_8474  <= TRANSPORT NOT a_SCOMMANDREG_F0_G  ;
and1_7457: n_8475 <=  gnd;
dff_7458: DFF_a8237

    PORT MAP ( D => a_EQ1177, CLK => a_STCSTATUS_F0_G_aCLK, CLRN => a_STCSTATUS_F0_G_aCLRN,
          PRN => vcc, Q => a_STCSTATUS_F0_G);
inv_7459: a_STCSTATUS_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7460: a_EQ1177 <=  n_8482  XOR n_8491;
or2_7461: n_8482 <=  n_8483  OR n_8487;
and3_7462: n_8483 <=  n_8484  AND n_8485  AND n_8486;
delay_7463: n_8484  <= TRANSPORT a_N2563_aNOT  ;
delay_7464: n_8485  <= TRANSPORT a_N2367  ;
delay_7465: n_8486  <= TRANSPORT a_N1530_aNOT  ;
and3_7466: n_8487 <=  n_8488  AND n_8489  AND n_8490;
delay_7467: n_8488  <= TRANSPORT a_N2563_aNOT  ;
inv_7468: n_8489  <= TRANSPORT NOT a_LC2_B15  ;
delay_7469: n_8490  <= TRANSPORT a_N1530_aNOT  ;
and1_7470: n_8491 <=  gnd;
delay_7471: n_8492  <= TRANSPORT clk  ;
filter_7472: FILTER_a8237

    PORT MAP (IN1 => n_8492, Y => a_STCSTATUS_F0_G_aCLK);
delay_7473: a_N1446  <= TRANSPORT a_EQ445  ;
xor2_7474: a_EQ445 <=  n_8496  XOR n_8503;
or2_7475: n_8496 <=  n_8497  OR n_8500;
and2_7476: n_8497 <=  n_8498  AND n_8499;
delay_7477: n_8498  <= TRANSPORT a_N57_aNOT  ;
delay_7478: n_8499  <= TRANSPORT a_N2565  ;
and2_7479: n_8500 <=  n_8501  AND n_8502;
delay_7480: n_8501  <= TRANSPORT a_N57_aNOT  ;
delay_7481: n_8502  <= TRANSPORT a_N2564  ;
and1_7482: n_8503 <=  gnd;
delay_7483: a_LC2_B22_aNOT  <= TRANSPORT a_EQ441  ;
xor2_7484: a_EQ441 <=  n_8506  XOR n_8516;
or2_7485: n_8506 <=  n_8507  OR n_8512;
and3_7486: n_8507 <=  n_8508  AND n_8509  AND n_8510;
delay_7487: n_8508  <= TRANSPORT a_N88_aNOT  ;
delay_7488: n_8509  <= TRANSPORT a_N1446  ;
delay_7489: n_8510  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
and3_7490: n_8512 <=  n_8513  AND n_8514  AND n_8515;
inv_7491: n_8513  <= TRANSPORT NOT a_N88_aNOT  ;
delay_7492: n_8514  <= TRANSPORT a_N1446  ;
delay_7493: n_8515  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and1_7494: n_8516 <=  gnd;
delay_7495: a_LC4_B19  <= TRANSPORT a_EQ539  ;
xor2_7496: a_EQ539 <=  n_8519  XOR n_8527;
or3_7497: n_8519 <=  n_8520  OR n_8522  OR n_8525;
and1_7498: n_8520 <=  n_8521;
delay_7499: n_8521  <= TRANSPORT a_LC2_B22_aNOT  ;
and2_7500: n_8522 <=  n_8523  AND n_8524;
delay_7501: n_8523  <= TRANSPORT a_N104_aNOT  ;
inv_7502: n_8524  <= TRANSPORT NOT dbin(1)  ;
and1_7503: n_8525 <=  n_8526;
delay_7504: n_8526  <= TRANSPORT a_N103_aNOT  ;
and1_7505: n_8527 <=  gnd;
delay_7506: a_LC1_B17  <= TRANSPORT a_LC1_B17_aIN  ;
xor2_7507: a_LC1_B17_aIN <=  n_8530  XOR n_8536;
or1_7508: n_8530 <=  n_8531;
and4_7509: n_8531 <=  n_8532  AND n_8533  AND n_8534  AND n_8535;
inv_7510: n_8532  <= TRANSPORT NOT a_N88_aNOT  ;
inv_7511: n_8533  <= TRANSPORT NOT a_N2564  ;
inv_7512: n_8534  <= TRANSPORT NOT a_N2565  ;
delay_7513: n_8535  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and1_7514: n_8536 <=  gnd;
delay_7515: a_LC2_B17_aNOT  <= TRANSPORT a_EQ444  ;
xor2_7516: a_EQ444 <=  n_8539  XOR n_8549;
or3_7517: n_8539 <=  n_8540  OR n_8543  OR n_8546;
and2_7518: n_8540 <=  n_8541  AND n_8542;
delay_7519: n_8541  <= TRANSPORT a_LC1_B17  ;
delay_7520: n_8542  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
and2_7521: n_8543 <=  n_8544  AND n_8545;
inv_7522: n_8544  <= TRANSPORT NOT a_N1119_aNOT  ;
delay_7523: n_8545  <= TRANSPORT a_LC1_B17  ;
and2_7524: n_8546 <=  n_8547  AND n_8548;
delay_7525: n_8547  <= TRANSPORT a_N57_aNOT  ;
delay_7526: n_8548  <= TRANSPORT a_LC1_B17  ;
and1_7527: n_8549 <=  gnd;
delay_7528: a_LC7_B17_aNOT  <= TRANSPORT a_EQ446  ;
xor2_7529: a_EQ446 <=  n_8552  XOR n_8561;
or2_7530: n_8552 <=  n_8553  OR n_8557;
and3_7531: n_8553 <=  n_8554  AND n_8555  AND n_8556;
inv_7532: n_8554  <= TRANSPORT NOT a_N57_aNOT  ;
inv_7533: n_8555  <= TRANSPORT NOT a_N84  ;
delay_7534: n_8556  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
and3_7535: n_8557 <=  n_8558  AND n_8559  AND n_8560;
inv_7536: n_8558  <= TRANSPORT NOT a_N2598_aNOT  ;
inv_7537: n_8559  <= TRANSPORT NOT a_N84  ;
delay_7538: n_8560  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
and1_7539: n_8561 <=  gnd;
delay_7540: a_LC6_B17_aNOT  <= TRANSPORT a_EQ440  ;
xor2_7541: a_EQ440 <=  n_8564  XOR n_8571;
or2_7542: n_8564 <=  n_8565  OR n_8567;
and1_7543: n_8565 <=  n_8566;
delay_7544: n_8566  <= TRANSPORT a_LC7_B17_aNOT  ;
and3_7545: n_8567 <=  n_8568  AND n_8569  AND n_8570;
inv_7546: n_8568  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7547: n_8569  <= TRANSPORT a_N84  ;
inv_7548: n_8570  <= TRANSPORT NOT dbin(2)  ;
and1_7549: n_8571 <=  gnd;
delay_7550: a_LC8_B17_aNOT  <= TRANSPORT a_EQ540  ;
xor2_7551: a_EQ540 <=  n_8574  XOR n_8582;
or3_7552: n_8574 <=  n_8575  OR n_8577  OR n_8579;
and1_7553: n_8575 <=  n_8576;
delay_7554: n_8576  <= TRANSPORT a_LC4_B19  ;
and1_7555: n_8577 <=  n_8578;
delay_7556: n_8578  <= TRANSPORT a_LC2_B17_aNOT  ;
and2_7557: n_8579 <=  n_8580  AND n_8581;
delay_7558: n_8580  <= TRANSPORT a_N2565  ;
delay_7559: n_8581  <= TRANSPORT a_LC6_B17_aNOT  ;
and1_7560: n_8582 <=  gnd;
delay_7561: a_N1432  <= TRANSPORT a_N1432_aIN  ;
xor2_7562: a_N1432_aIN <=  n_8585  XOR n_8589;
or1_7563: n_8585 <=  n_8586;
and2_7564: n_8586 <=  n_8587  AND n_8588;
delay_7565: n_8587  <= TRANSPORT a_N2563_aNOT  ;
delay_7566: n_8588  <= TRANSPORT a_N1119_aNOT  ;
and1_7567: n_8589 <=  gnd;
delay_7568: a_N1442_aNOT  <= TRANSPORT a_EQ442  ;
xor2_7569: a_EQ442 <=  n_8592  XOR n_8601;
or2_7570: n_8592 <=  n_8593  OR n_8597;
and3_7571: n_8593 <=  n_8594  AND n_8595  AND n_8596;
inv_7572: n_8594  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7573: n_8595  <= TRANSPORT a_N1432  ;
delay_7574: n_8596  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
and3_7575: n_8597 <=  n_8598  AND n_8599  AND n_8600;
delay_7576: n_8598  <= TRANSPORT a_N88_aNOT  ;
delay_7577: n_8599  <= TRANSPORT a_N1432  ;
delay_7578: n_8600  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
and1_7579: n_8601 <=  gnd;
dff_7580: DFF_a8237

    PORT MAP ( D => a_EQ1158, CLK => a_SMASKREG_F1_G_aNOT_aCLK, CLRN => a_SMASKREG_F1_G_aNOT_aCLRN,
          PRN => vcc, Q => a_SMASKREG_F1_G_aNOT);
inv_7581: a_SMASKREG_F1_G_aNOT_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7582: a_EQ1158 <=  n_8608  XOR n_8614;
or2_7583: n_8608 <=  n_8609  OR n_8612;
and2_7584: n_8609 <=  n_8610  AND n_8611;
delay_7585: n_8610  <= TRANSPORT a_N2563_aNOT  ;
delay_7586: n_8611  <= TRANSPORT a_LC8_B17_aNOT  ;
and1_7587: n_8612 <=  n_8613;
delay_7588: n_8613  <= TRANSPORT a_N1442_aNOT  ;
and1_7589: n_8614 <=  gnd;
delay_7590: n_8615  <= TRANSPORT clk  ;
filter_7591: FILTER_a8237

    PORT MAP (IN1 => n_8615, Y => a_SMASKREG_F1_G_aNOT_aCLK);
delay_7592: a_LC4_B9_aNOT  <= TRANSPORT a_LC4_B9_aNOT_aIN  ;
xor2_7593: a_LC4_B9_aNOT_aIN <=  n_8619  XOR n_8625;
or1_7594: n_8619 <=  n_8620;
and4_7595: n_8620 <=  n_8621  AND n_8622  AND n_8623  AND n_8624;
inv_7596: n_8621  <= TRANSPORT NOT a_N87  ;
inv_7597: n_8622  <= TRANSPORT NOT a_N63_aNOT  ;
inv_7598: n_8623  <= TRANSPORT NOT dbin(0)  ;
delay_7599: n_8624  <= TRANSPORT dbin(1)  ;
and1_7600: n_8625 <=  gnd;
dff_7601: DFF_a8237

    PORT MAP ( D => a_EQ1175, CLK => a_SREQUESTREG_F2_G_aCLK, CLRN => a_SREQUESTREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SREQUESTREG_F2_G);
inv_7602: a_SREQUESTREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7603: a_EQ1175 <=  n_8633  XOR n_8642;
or2_7604: n_8633 <=  n_8634  OR n_8638;
and3_7605: n_8634 <=  n_8635  AND n_8636  AND n_8637;
delay_7606: n_8635  <= TRANSPORT a_N2563_aNOT  ;
delay_7607: n_8636  <= TRANSPORT a_LC4_B9_aNOT  ;
delay_7608: n_8637  <= TRANSPORT dbin(2)  ;
and3_7609: n_8638 <=  n_8639  AND n_8640  AND n_8641;
delay_7610: n_8639  <= TRANSPORT a_N2563_aNOT  ;
inv_7611: n_8640  <= TRANSPORT NOT a_LC4_B9_aNOT  ;
delay_7612: n_8641  <= TRANSPORT a_SREQUESTREG_F2_G  ;
and1_7613: n_8642 <=  gnd;
delay_7614: n_8643  <= TRANSPORT clk  ;
filter_7615: FILTER_a8237

    PORT MAP (IN1 => n_8643, Y => a_SREQUESTREG_F2_G_aCLK);
dff_7616: DFF_a8237

    PORT MAP ( D => a_EQ1179, CLK => a_STCSTATUS_F2_G_aCLK, CLRN => a_STCSTATUS_F2_G_aCLRN,
          PRN => vcc, Q => a_STCSTATUS_F2_G);
inv_7617: a_STCSTATUS_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7618: a_EQ1179 <=  n_8652  XOR n_8660;
or2_7619: n_8652 <=  n_8653  OR n_8656;
and2_7620: n_8653 <=  n_8654  AND n_8655;
delay_7621: n_8654  <= TRANSPORT a_N2592  ;
delay_7622: n_8655  <= TRANSPORT a_STCSTATUS_F2_G  ;
and3_7623: n_8656 <=  n_8657  AND n_8658  AND n_8659;
inv_7624: n_8657  <= TRANSPORT NOT a_N2376  ;
delay_7625: n_8658  <= TRANSPORT a_N57_aNOT  ;
delay_7626: n_8659  <= TRANSPORT a_N2592  ;
and1_7627: n_8660 <=  gnd;
delay_7628: n_8661  <= TRANSPORT clk  ;
filter_7629: FILTER_a8237

    PORT MAP (IN1 => n_8661, Y => a_STCSTATUS_F2_G_aCLK);
delay_7630: a_LC3_B19_aNOT  <= TRANSPORT a_LC3_B19_aNOT_aIN  ;
xor2_7631: a_LC3_B19_aNOT_aIN <=  n_8665  XOR n_8671;
or1_7632: n_8665 <=  n_8666;
and4_7633: n_8666 <=  n_8667  AND n_8668  AND n_8669  AND n_8670;
inv_7634: n_8667  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7635: n_8668  <= TRANSPORT a_N2565  ;
inv_7636: n_8669  <= TRANSPORT NOT dbin(0)  ;
delay_7637: n_8670  <= TRANSPORT dbin(1)  ;
and1_7638: n_8671 <=  gnd;
delay_7639: a_LC7_B19  <= TRANSPORT a_EQ536  ;
xor2_7640: a_EQ536 <=  n_8674  XOR n_8683;
or3_7641: n_8674 <=  n_8675  OR n_8678  OR n_8681;
and2_7642: n_8675 <=  n_8676  AND n_8677;
inv_7643: n_8676  <= TRANSPORT NOT dbin(2)  ;
delay_7644: n_8677  <= TRANSPORT a_LC3_B19_aNOT  ;
and2_7645: n_8678 <=  n_8679  AND n_8680;
delay_7646: n_8679  <= TRANSPORT a_N104_aNOT  ;
inv_7647: n_8680  <= TRANSPORT NOT dbin(2)  ;
and1_7648: n_8681 <=  n_8682;
delay_7649: n_8682  <= TRANSPORT a_N103_aNOT  ;
and1_7650: n_8683 <=  gnd;
delay_7651: a_LC2_B19  <= TRANSPORT a_EQ435  ;
xor2_7652: a_EQ435 <=  n_8686  XOR n_8696;
or2_7653: n_8686 <=  n_8687  OR n_8692;
and3_7654: n_8687 <=  n_8688  AND n_8689  AND n_8690;
delay_7655: n_8688  <= TRANSPORT a_N2565  ;
inv_7656: n_8689  <= TRANSPORT NOT dbin(1)  ;
delay_7657: n_8690  <= TRANSPORT a_SMASKREG_F2_G_aNOT  ;
and3_7658: n_8692 <=  n_8693  AND n_8694  AND n_8695;
delay_7659: n_8693  <= TRANSPORT a_N2565  ;
delay_7660: n_8694  <= TRANSPORT dbin(0)  ;
delay_7661: n_8695  <= TRANSPORT a_SMASKREG_F2_G_aNOT  ;
and1_7662: n_8696 <=  gnd;
delay_7663: a_LC6_B19  <= TRANSPORT a_EQ537  ;
xor2_7664: a_EQ537 <=  n_8699  XOR n_8708;
or3_7665: n_8699 <=  n_8700  OR n_8702  OR n_8705;
and1_7666: n_8700 <=  n_8701;
delay_7667: n_8701  <= TRANSPORT a_LC7_B19  ;
and2_7668: n_8702 <=  n_8703  AND n_8704;
delay_7669: n_8703  <= TRANSPORT a_LC2_B19  ;
inv_7670: n_8704  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and2_7671: n_8705 <=  n_8706  AND n_8707;
inv_7672: n_8706  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7673: n_8707  <= TRANSPORT a_LC2_B19  ;
and1_7674: n_8708 <=  gnd;
delay_7675: a_N46  <= TRANSPORT a_N46_aIN  ;
xor2_7676: a_N46_aIN <=  n_8711  XOR n_8715;
or1_7677: n_8711 <=  n_8712;
and2_7678: n_8712 <=  n_8713  AND n_8714;
inv_7679: n_8713  <= TRANSPORT NOT a_N2564  ;
inv_7680: n_8714  <= TRANSPORT NOT a_N2565  ;
and1_7681: n_8715 <=  gnd;
delay_7682: a_LC6_B22_aNOT  <= TRANSPORT a_EQ535  ;
xor2_7683: a_EQ535 <=  n_8718  XOR n_8728;
or3_7684: n_8718 <=  n_8719  OR n_8722  OR n_8725;
and2_7685: n_8719 <=  n_8720  AND n_8721;
inv_7686: n_8720  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7687: n_8721  <= TRANSPORT a_N46  ;
and2_7688: n_8722 <=  n_8723  AND n_8724;
delay_7689: n_8723  <= TRANSPORT a_N57_aNOT  ;
inv_7690: n_8724  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and2_7691: n_8725 <=  n_8726  AND n_8727;
delay_7692: n_8726  <= TRANSPORT a_N57_aNOT  ;
delay_7693: n_8727  <= TRANSPORT a_SCHANNEL_F0_G  ;
and1_7694: n_8728 <=  gnd;
delay_7695: a_LC5_B22_aNOT  <= TRANSPORT a_EQ538  ;
xor2_7696: a_EQ538 <=  n_8731  XOR n_8739;
or2_7697: n_8731 <=  n_8732  OR n_8735;
and2_7698: n_8732 <=  n_8733  AND n_8734;
delay_7699: n_8733  <= TRANSPORT a_N2563_aNOT  ;
delay_7700: n_8734  <= TRANSPORT a_LC6_B19  ;
and3_7701: n_8735 <=  n_8736  AND n_8737  AND n_8738;
delay_7702: n_8736  <= TRANSPORT a_N2563_aNOT  ;
delay_7703: n_8737  <= TRANSPORT a_LC6_B22_aNOT  ;
delay_7704: n_8738  <= TRANSPORT a_SMASKREG_F2_G_aNOT  ;
and1_7705: n_8739 <=  gnd;
delay_7706: a_LC8_B22_aNOT  <= TRANSPORT a_EQ436  ;
xor2_7707: a_EQ436 <=  n_8742  XOR n_8751;
or2_7708: n_8742 <=  n_8743  OR n_8747;
and3_7709: n_8743 <=  n_8744  AND n_8745  AND n_8746;
delay_7710: n_8744  <= TRANSPORT a_N2563_aNOT  ;
delay_7711: n_8745  <= TRANSPORT a_N1119_aNOT  ;
delay_7712: n_8746  <= TRANSPORT a_SMASKREG_F2_G_aNOT  ;
and3_7713: n_8747 <=  n_8748  AND n_8749  AND n_8750;
delay_7714: n_8748  <= TRANSPORT a_N2563_aNOT  ;
delay_7715: n_8749  <= TRANSPORT a_N57_aNOT  ;
delay_7716: n_8750  <= TRANSPORT a_N1119_aNOT  ;
and1_7717: n_8751 <=  gnd;
delay_7718: a_LC7_B22_aNOT  <= TRANSPORT a_EQ534  ;
xor2_7719: a_EQ534 <=  n_8754  XOR n_8761;
or2_7720: n_8754 <=  n_8755  OR n_8757;
and1_7721: n_8755 <=  n_8756;
delay_7722: n_8756  <= TRANSPORT a_LC8_B22_aNOT  ;
and3_7723: n_8757 <=  n_8758  AND n_8759  AND n_8760;
delay_7724: n_8758  <= TRANSPORT a_N2563_aNOT  ;
delay_7725: n_8759  <= TRANSPORT a_N2377  ;
delay_7726: n_8760  <= TRANSPORT a_N1446  ;
and1_7727: n_8761 <=  gnd;
dff_7728: DFF_a8237

    PORT MAP ( D => a_EQ1159, CLK => a_SMASKREG_F2_G_aNOT_aCLK, CLRN => a_SMASKREG_F2_G_aNOT_aCLRN,
          PRN => vcc, Q => a_SMASKREG_F2_G_aNOT);
inv_7729: a_SMASKREG_F2_G_aNOT_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7730: a_EQ1159 <=  n_8768  XOR n_8775;
or2_7731: n_8768 <=  n_8769  OR n_8771;
and1_7732: n_8769 <=  n_8770;
delay_7733: n_8770  <= TRANSPORT a_LC5_B22_aNOT  ;
and3_7734: n_8771 <=  n_8772  AND n_8773  AND n_8774;
inv_7735: n_8772  <= TRANSPORT NOT a_N2376  ;
delay_7736: n_8773  <= TRANSPORT a_LC7_B22_aNOT  ;
delay_7737: n_8774  <= TRANSPORT a_SCH2MODEREG_F2_G  ;
and1_7738: n_8775 <=  gnd;
delay_7739: n_8776  <= TRANSPORT clk  ;
filter_7740: FILTER_a8237

    PORT MAP (IN1 => n_8776, Y => a_SMASKREG_F2_G_aNOT_aCLK);
delay_7741: a_N2571_aNOT  <= TRANSPORT a_EQ624  ;
xor2_7742: a_EQ624 <=  n_8780  XOR n_8785;
or2_7743: n_8780 <=  n_8781  OR n_8783;
and1_7744: n_8781 <=  n_8782;
delay_7745: n_8782  <= TRANSPORT a_N2367  ;
and1_7746: n_8783 <=  n_8784;
delay_7747: n_8784  <= TRANSPORT a_N87  ;
and1_7748: n_8785 <=  gnd;
dff_7749: DFF_a8237

    PORT MAP ( D => a_EQ1125, CLK => a_SCOMMANDREG_F2_G_aCLK, CLRN => a_SCOMMANDREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F2_G);
inv_7750: a_SCOMMANDREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7751: a_EQ1125 <=  n_8793  XOR n_8801;
or2_7752: n_8793 <=  n_8794  OR n_8798;
and3_7753: n_8794 <=  n_8795  AND n_8796  AND n_8797;
delay_7754: n_8795  <= TRANSPORT a_N2563_aNOT  ;
delay_7755: n_8796  <= TRANSPORT a_N2571_aNOT  ;
delay_7756: n_8797  <= TRANSPORT a_SCOMMANDREG_F2_G  ;
and2_7757: n_8798 <=  n_8799  AND n_8800;
delay_7758: n_8799  <= TRANSPORT dbin(2)  ;
inv_7759: n_8800  <= TRANSPORT NOT a_N2571_aNOT  ;
and1_7760: n_8801 <=  gnd;
delay_7761: n_8802  <= TRANSPORT clk  ;
filter_7762: FILTER_a8237

    PORT MAP (IN1 => n_8802, Y => a_SCOMMANDREG_F2_G_aCLK);
delay_7763: a_LC5_B8_aNOT  <= TRANSPORT a_EQ466  ;
xor2_7764: a_EQ466 <=  n_8806  XOR n_8812;
or2_7765: n_8806 <=  n_8807  OR n_8809;
and1_7766: n_8807 <=  n_8808;
inv_7767: n_8808  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and2_7768: n_8809 <=  n_8810  AND n_8811;
delay_7769: n_8810  <= TRANSPORT a_N2377  ;
delay_7770: n_8811  <= TRANSPORT a_SCH3MODEREG_F2_G  ;
and1_7771: n_8812 <=  gnd;
delay_7772: a_N1565  <= TRANSPORT a_EQ464  ;
xor2_7773: a_EQ464 <=  n_8815  XOR n_8824;
or4_7774: n_8815 <=  n_8816  OR n_8818  OR n_8820  OR n_8822;
and1_7775: n_8816 <=  n_8817;
inv_7776: n_8817  <= TRANSPORT NOT dbin(1)  ;
and1_7777: n_8818 <=  n_8819;
inv_7778: n_8819  <= TRANSPORT NOT dbin(0)  ;
and1_7779: n_8820 <=  n_8821;
inv_7780: n_8821  <= TRANSPORT NOT dbin(2)  ;
and1_7781: n_8822 <=  n_8823;
inv_7782: n_8823  <= TRANSPORT NOT a_N2565  ;
and1_7783: n_8824 <=  gnd;
delay_7784: a_LC4_B8  <= TRANSPORT a_EQ467  ;
xor2_7785: a_EQ467 <=  n_8827  XOR n_8835;
or2_7786: n_8827 <=  n_8828  OR n_8831;
and2_7787: n_8828 <=  n_8829  AND n_8830;
delay_7788: n_8829  <= TRANSPORT a_N57_aNOT  ;
delay_7789: n_8830  <= TRANSPORT a_LC5_B8_aNOT  ;
and3_7790: n_8831 <=  n_8832  AND n_8833  AND n_8834;
inv_7791: n_8832  <= TRANSPORT NOT a_N57_aNOT  ;
inv_7792: n_8833  <= TRANSPORT NOT a_N2564  ;
delay_7793: n_8834  <= TRANSPORT a_N1565  ;
and1_7794: n_8835 <=  gnd;
delay_7795: a_N1563_aNOT  <= TRANSPORT a_EQ463  ;
xor2_7796: a_EQ463 <=  n_8838  XOR n_8847;
or2_7797: n_8838 <=  n_8839  OR n_8843;
and2_7798: n_8839 <=  n_8840  AND n_8841;
delay_7799: n_8840  <= TRANSPORT a_LC4_B8  ;
delay_7800: n_8841  <= TRANSPORT a_SMASKREG_F3_G_aNOT  ;
and3_7801: n_8843 <=  n_8844  AND n_8845  AND n_8846;
inv_7802: n_8844  <= TRANSPORT NOT a_N2376  ;
delay_7803: n_8845  <= TRANSPORT a_N57_aNOT  ;
delay_7804: n_8846  <= TRANSPORT a_SMASKREG_F3_G_aNOT  ;
and1_7805: n_8847 <=  gnd;
delay_7806: a_N24  <= TRANSPORT a_EQ177  ;
xor2_7807: a_EQ177 <=  n_8850  XOR n_8857;
or3_7808: n_8850 <=  n_8851  OR n_8853  OR n_8855;
and1_7809: n_8851 <=  n_8852;
inv_7810: n_8852  <= TRANSPORT NOT dbin(1)  ;
and1_7811: n_8853 <=  n_8854;
inv_7812: n_8854  <= TRANSPORT NOT dbin(0)  ;
and1_7813: n_8855 <=  n_8856;
delay_7814: n_8856  <= TRANSPORT dbin(2)  ;
and1_7815: n_8857 <=  gnd;
delay_7816: a_LC2_B8_aNOT  <= TRANSPORT a_EQ461  ;
xor2_7817: a_EQ461 <=  n_8860  XOR n_8867;
or2_7818: n_8860 <=  n_8861  OR n_8864;
and2_7819: n_8861 <=  n_8862  AND n_8863;
delay_7820: n_8862  <= TRANSPORT a_N2565  ;
inv_7821: n_8863  <= TRANSPORT NOT a_N24  ;
and2_7822: n_8864 <=  n_8865  AND n_8866;
delay_7823: n_8865  <= TRANSPORT a_N2564  ;
inv_7824: n_8866  <= TRANSPORT NOT dbin(3)  ;
and1_7825: n_8867 <=  gnd;
delay_7826: a_LC1_B8  <= TRANSPORT a_EQ462  ;
xor2_7827: a_EQ462 <=  n_8870  XOR n_8878;
or3_7828: n_8870 <=  n_8871  OR n_8873  OR n_8876;
and1_7829: n_8871 <=  n_8872;
delay_7830: n_8872  <= TRANSPORT a_N1563_aNOT  ;
and2_7831: n_8873 <=  n_8874  AND n_8875;
inv_7832: n_8874  <= TRANSPORT NOT a_N57_aNOT  ;
delay_7833: n_8875  <= TRANSPORT a_LC2_B8_aNOT  ;
and1_7834: n_8876 <=  n_8877;
delay_7835: n_8877  <= TRANSPORT a_N103_aNOT  ;
and1_7836: n_8878 <=  gnd;
dff_7837: DFF_a8237

    PORT MAP ( D => a_EQ1160, CLK => a_SMASKREG_F3_G_aNOT_aCLK, CLRN => a_SMASKREG_F3_G_aNOT_aCLRN,
          PRN => vcc, Q => a_SMASKREG_F3_G_aNOT);
inv_7838: a_SMASKREG_F3_G_aNOT_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7839: a_EQ1160 <=  n_8885  XOR n_8893;
or2_7840: n_8885 <=  n_8886  OR n_8889;
and2_7841: n_8886 <=  n_8887  AND n_8888;
delay_7842: n_8887  <= TRANSPORT a_N2563_aNOT  ;
delay_7843: n_8888  <= TRANSPORT a_LC1_B8  ;
and3_7844: n_8889 <=  n_8890  AND n_8891  AND n_8892;
delay_7845: n_8890  <= TRANSPORT a_N2563_aNOT  ;
inv_7846: n_8891  <= TRANSPORT NOT a_N2377  ;
delay_7847: n_8892  <= TRANSPORT a_N2528  ;
and1_7848: n_8893 <=  gnd;
delay_7849: n_8894  <= TRANSPORT clk  ;
filter_7850: FILTER_a8237

    PORT MAP (IN1 => n_8894, Y => a_SMASKREG_F3_G_aNOT_aCLK);
dff_7851: DFF_a8237

    PORT MAP ( D => a_EQ1180, CLK => a_STCSTATUS_F3_G_aCLK, CLRN => a_STCSTATUS_F3_G_aCLRN,
          PRN => vcc, Q => a_STCSTATUS_F3_G);
inv_7852: a_STCSTATUS_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7853: a_EQ1180 <=  n_8903  XOR n_8911;
or2_7854: n_8903 <=  n_8904  OR n_8907;
and2_7855: n_8904 <=  n_8905  AND n_8906;
delay_7856: n_8905  <= TRANSPORT a_N2592  ;
delay_7857: n_8906  <= TRANSPORT a_STCSTATUS_F3_G  ;
and3_7858: n_8907 <=  n_8908  AND n_8909  AND n_8910;
inv_7859: n_8908  <= TRANSPORT NOT a_N2377  ;
delay_7860: n_8909  <= TRANSPORT a_N57_aNOT  ;
delay_7861: n_8910  <= TRANSPORT a_N2592  ;
and1_7862: n_8911 <=  gnd;
delay_7863: n_8912  <= TRANSPORT clk  ;
filter_7864: FILTER_a8237

    PORT MAP (IN1 => n_8912, Y => a_STCSTATUS_F3_G_aCLK);
delay_7865: a_LC3_B18  <= TRANSPORT a_EQ541  ;
xor2_7866: a_EQ541 <=  n_8916  XOR n_8924;
or2_7867: n_8916 <=  n_8917  OR n_8920;
and1_7868: n_8917 <=  n_8918;
delay_7869: n_8918  <= TRANSPORT a_SREQUESTREG_F3_G  ;
and3_7870: n_8920 <=  n_8921  AND n_8922  AND n_8923;
inv_7871: n_8921  <= TRANSPORT NOT a_N2566_aNOT  ;
delay_7872: n_8922  <= TRANSPORT dbin(0)  ;
delay_7873: n_8923  <= TRANSPORT dbin(1)  ;
and1_7874: n_8924 <=  gnd;
dff_7875: DFF_a8237

    PORT MAP ( D => a_EQ1176, CLK => a_SREQUESTREG_F3_G_aCLK, CLRN => a_SREQUESTREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SREQUESTREG_F3_G);
inv_7876: a_SREQUESTREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7877: a_EQ1176 <=  n_8931  XOR n_8940;
or2_7878: n_8931 <=  n_8932  OR n_8936;
and3_7879: n_8932 <=  n_8933  AND n_8934  AND n_8935;
delay_7880: n_8933  <= TRANSPORT a_N2563_aNOT  ;
delay_7881: n_8934  <= TRANSPORT a_N24  ;
delay_7882: n_8935  <= TRANSPORT a_LC3_B18  ;
and3_7883: n_8936 <=  n_8937  AND n_8938  AND n_8939;
delay_7884: n_8937  <= TRANSPORT a_N2563_aNOT  ;
delay_7885: n_8938  <= TRANSPORT a_N2566_aNOT  ;
delay_7886: n_8939  <= TRANSPORT a_LC3_B18  ;
and1_7887: n_8940 <=  gnd;
delay_7888: n_8941  <= TRANSPORT clk  ;
filter_7889: FILTER_a8237

    PORT MAP (IN1 => n_8941, Y => a_SREQUESTREG_F3_G_aCLK);
dff_7890: DFF_a8237

    PORT MAP ( D => a_EQ1126, CLK => a_SCOMMANDREG_F3_G_aCLK, CLRN => a_SCOMMANDREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F3_G);
inv_7891: a_SCOMMANDREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7892: a_EQ1126 <=  n_8950  XOR n_8958;
or2_7893: n_8950 <=  n_8951  OR n_8955;
and3_7894: n_8951 <=  n_8952  AND n_8953  AND n_8954;
delay_7895: n_8952  <= TRANSPORT a_N2563_aNOT  ;
delay_7896: n_8953  <= TRANSPORT a_N2571_aNOT  ;
delay_7897: n_8954  <= TRANSPORT a_SCOMMANDREG_F3_G  ;
and2_7898: n_8955 <=  n_8956  AND n_8957;
inv_7899: n_8956  <= TRANSPORT NOT a_N2571_aNOT  ;
delay_7900: n_8957  <= TRANSPORT dbin(3)  ;
and1_7901: n_8958 <=  gnd;
delay_7902: n_8959  <= TRANSPORT clk  ;
filter_7903: FILTER_a8237

    PORT MAP (IN1 => n_8959, Y => a_SCOMMANDREG_F3_G_aCLK);
dff_7904: DFF_a8237

    PORT MAP ( D => a_EQ1127, CLK => a_SCOMMANDREG_F4_G_aCLK, CLRN => a_SCOMMANDREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F4_G);
inv_7905: a_SCOMMANDREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7906: a_EQ1127 <=  n_8968  XOR n_8976;
or2_7907: n_8968 <=  n_8969  OR n_8973;
and3_7908: n_8969 <=  n_8970  AND n_8971  AND n_8972;
delay_7909: n_8970  <= TRANSPORT a_N2563_aNOT  ;
delay_7910: n_8971  <= TRANSPORT a_N2571_aNOT  ;
delay_7911: n_8972  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
and2_7912: n_8973 <=  n_8974  AND n_8975;
inv_7913: n_8974  <= TRANSPORT NOT a_N2571_aNOT  ;
delay_7914: n_8975  <= TRANSPORT dbin(4)  ;
and1_7915: n_8976 <=  gnd;
delay_7916: n_8977  <= TRANSPORT clk  ;
filter_7917: FILTER_a8237

    PORT MAP (IN1 => n_8977, Y => a_SCOMMANDREG_F4_G_aCLK);
dff_7918: DFF_a8237

    PORT MAP ( D => a_EQ1112, CLK => a_SCH3MODEREG_F5_G_aCLK, CLRN => a_SCH3MODEREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH3MODEREG_F5_G);
inv_7919: a_SCH3MODEREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7920: a_EQ1112 <=  n_8986  XOR n_8993;
or2_7921: n_8986 <=  n_8987  OR n_8990;
and2_7922: n_8987 <=  n_8988  AND n_8989;
inv_7923: n_8988  <= TRANSPORT NOT a_N2570_aNOT  ;
delay_7924: n_8989  <= TRANSPORT dbin(7)  ;
and2_7925: n_8990 <=  n_8991  AND n_8992;
delay_7926: n_8991  <= TRANSPORT a_N2570_aNOT  ;
delay_7927: n_8992  <= TRANSPORT a_SCH3MODEREG_F5_G  ;
and1_7928: n_8993 <=  gnd;
delay_7929: n_8994  <= TRANSPORT clk  ;
filter_7930: FILTER_a8237

    PORT MAP (IN1 => n_8994, Y => a_SCH3MODEREG_F5_G_aCLK);
dff_7931: DFF_a8237

    PORT MAP ( D => a_EQ984, CLK => a_SCH1MODEREG_F5_G_aCLK, CLRN => a_SCH1MODEREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH1MODEREG_F5_G);
inv_7932: a_SCH1MODEREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7933: a_EQ984 <=  n_9003  XOR n_9010;
or2_7934: n_9003 <=  n_9004  OR n_9007;
and2_7935: n_9004 <=  n_9005  AND n_9006;
inv_7936: n_9005  <= TRANSPORT NOT a_N2568  ;
delay_7937: n_9006  <= TRANSPORT a_SCH1MODEREG_F5_G  ;
and2_7938: n_9007 <=  n_9008  AND n_9009;
delay_7939: n_9008  <= TRANSPORT a_N2568  ;
delay_7940: n_9009  <= TRANSPORT dbin(7)  ;
and1_7941: n_9010 <=  gnd;
delay_7942: n_9011  <= TRANSPORT clk  ;
filter_7943: FILTER_a8237

    PORT MAP (IN1 => n_9011, Y => a_SCH1MODEREG_F5_G_aCLK);
dff_7944: DFF_a8237

    PORT MAP ( D => a_EQ1048, CLK => a_SCH2MODEREG_F5_G_aCLK, CLRN => a_SCH2MODEREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH2MODEREG_F5_G);
inv_7945: a_SCH2MODEREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7946: a_EQ1048 <=  n_9020  XOR n_9027;
or2_7947: n_9020 <=  n_9021  OR n_9024;
and2_7948: n_9021 <=  n_9022  AND n_9023;
inv_7949: n_9022  <= TRANSPORT NOT a_N2569_aNOT  ;
delay_7950: n_9023  <= TRANSPORT dbin(7)  ;
and2_7951: n_9024 <=  n_9025  AND n_9026;
delay_7952: n_9025  <= TRANSPORT a_N2569_aNOT  ;
delay_7953: n_9026  <= TRANSPORT a_SCH2MODEREG_F5_G  ;
and1_7954: n_9027 <=  gnd;
delay_7955: n_9028  <= TRANSPORT clk  ;
filter_7956: FILTER_a8237

    PORT MAP (IN1 => n_9028, Y => a_SCH2MODEREG_F5_G_aCLK);
delay_7957: a_LC1_B15  <= TRANSPORT a_EQ533  ;
xor2_7958: a_EQ533 <=  n_9032  XOR n_9042;
or3_7959: n_9032 <=  n_9033  OR n_9036  OR n_9039;
and2_7960: n_9033 <=  n_9034  AND n_9035;
delay_7961: n_9034  <= TRANSPORT a_N2563_aNOT  ;
delay_7962: n_9035  <= TRANSPORT a_N75_aNOT  ;
and2_7963: n_9036 <=  n_9037  AND n_9038;
delay_7964: n_9037  <= TRANSPORT a_N2563_aNOT  ;
delay_7965: n_9038  <= TRANSPORT ncs  ;
and2_7966: n_9039 <=  n_9040  AND n_9041;
delay_7967: n_9040  <= TRANSPORT a_N2563_aNOT  ;
delay_7968: n_9041  <= TRANSPORT niorin  ;
and1_7969: n_9042 <=  gnd;
delay_7970: a_N2390  <= TRANSPORT a_N2390_aIN  ;
xor2_7971: a_N2390_aIN <=  n_9045  XOR n_9049;
or1_7972: n_9045 <=  n_9046;
and2_7973: n_9046 <=  n_9047  AND n_9048;
delay_7974: n_9047  <= TRANSPORT a_LC2_B15  ;
delay_7975: n_9048  <= TRANSPORT a_N66  ;
and1_7976: n_9049 <=  gnd;
dff_7977: DFF_a8237

    PORT MAP ( D => a_EQ1162, CLK => a_SMODECOUNTER_F1_G_aCLK, CLRN => a_SMODECOUNTER_F1_G_aCLRN,
          PRN => vcc, Q => a_SMODECOUNTER_F1_G);
inv_7978: a_SMODECOUNTER_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7979: a_EQ1162 <=  n_9057  XOR n_9072;
or3_7980: n_9057 <=  n_9058  OR n_9063  OR n_9067;
and3_7981: n_9058 <=  n_9059  AND n_9060  AND n_9061;
delay_7982: n_9059  <= TRANSPORT a_LC1_B15  ;
delay_7983: n_9060  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_7984: n_9061  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and3_7985: n_9063 <=  n_9064  AND n_9065  AND n_9066;
delay_7986: n_9064  <= TRANSPORT a_LC1_B15  ;
inv_7987: n_9065  <= TRANSPORT NOT a_N2390  ;
delay_7988: n_9066  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
and4_7989: n_9067 <=  n_9068  AND n_9069  AND n_9070  AND n_9071;
delay_7990: n_9068  <= TRANSPORT a_LC1_B15  ;
delay_7991: n_9069  <= TRANSPORT a_N2390  ;
inv_7992: n_9070  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_7993: n_9071  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and1_7994: n_9072 <=  gnd;
delay_7995: n_9073  <= TRANSPORT clk  ;
filter_7996: FILTER_a8237

    PORT MAP (IN1 => n_9073, Y => a_SMODECOUNTER_F1_G_aCLK);
dff_7997: DFF_a8237

    PORT MAP ( D => a_EQ1161, CLK => a_SMODECOUNTER_F0_G_aCLK, CLRN => a_SMODECOUNTER_F0_G_aCLRN,
          PRN => vcc, Q => a_SMODECOUNTER_F0_G);
inv_7998: a_SMODECOUNTER_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_7999: a_EQ1161 <=  n_9081  XOR n_9095;
or3_8000: n_9081 <=  n_9082  OR n_9086  OR n_9090;
and3_8001: n_9082 <=  n_9083  AND n_9084  AND n_9085;
inv_8002: n_9083  <= TRANSPORT NOT a_LC2_B15  ;
delay_8003: n_9084  <= TRANSPORT a_LC1_B15  ;
delay_8004: n_9085  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and3_8005: n_9086 <=  n_9087  AND n_9088  AND n_9089;
inv_8006: n_9087  <= TRANSPORT NOT a_N66  ;
delay_8007: n_9088  <= TRANSPORT a_LC1_B15  ;
delay_8008: n_9089  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and4_8009: n_9090 <=  n_9091  AND n_9092  AND n_9093  AND n_9094;
delay_8010: n_9091  <= TRANSPORT a_LC2_B15  ;
delay_8011: n_9092  <= TRANSPORT a_N66  ;
delay_8012: n_9093  <= TRANSPORT a_LC1_B15  ;
inv_8013: n_9094  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and1_8014: n_9095 <=  gnd;
delay_8015: n_9096  <= TRANSPORT clk  ;
filter_8016: FILTER_a8237

    PORT MAP (IN1 => n_9096, Y => a_SMODECOUNTER_F0_G_aCLK);
dff_8017: DFF_a8237

    PORT MAP ( D => a_EQ920, CLK => a_SCH0MODEREG_F5_G_aCLK, CLRN => a_SCH0MODEREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH0MODEREG_F5_G);
inv_8018: a_SCH0MODEREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8019: a_EQ920 <=  n_9105  XOR n_9112;
or2_8020: n_9105 <=  n_9106  OR n_9109;
and2_8021: n_9106 <=  n_9107  AND n_9108;
inv_8022: n_9107  <= TRANSPORT NOT a_N2567  ;
delay_8023: n_9108  <= TRANSPORT a_SCH0MODEREG_F5_G  ;
and2_8024: n_9109 <=  n_9110  AND n_9111;
delay_8025: n_9110  <= TRANSPORT a_N2567  ;
delay_8026: n_9111  <= TRANSPORT dbin(7)  ;
and1_8027: n_9112 <=  gnd;
delay_8028: n_9113  <= TRANSPORT clk  ;
filter_8029: FILTER_a8237

    PORT MAP (IN1 => n_9113, Y => a_SCH0MODEREG_F5_G_aCLK);
dff_8030: DFF_a8237

    PORT MAP ( D => a_EQ1011, CLK => a_SCH2BAROUT_F0_G_aCLK, CLRN => a_SCH2BAROUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F0_G);
inv_8031: a_SCH2BAROUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8032: a_EQ1011 <=  n_9122  XOR n_9129;
or2_8033: n_9122 <=  n_9123  OR n_9126;
and2_8034: n_9123 <=  n_9124  AND n_9125;
delay_8035: n_9124  <= TRANSPORT a_N2582_aNOT  ;
delay_8036: n_9125  <= TRANSPORT a_SCH2BAROUT_F0_G  ;
and2_8037: n_9126 <=  n_9127  AND n_9128;
inv_8038: n_9127  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8039: n_9128  <= TRANSPORT dbin(0)  ;
and1_8040: n_9129 <=  gnd;
delay_8041: n_9130  <= TRANSPORT clk  ;
filter_8042: FILTER_a8237

    PORT MAP (IN1 => n_9130, Y => a_SCH2BAROUT_F0_G_aCLK);
dff_8043: DFF_a8237

    PORT MAP ( D => a_EQ1045, CLK => a_SCH2MODEREG_F2_G_aCLK, CLRN => a_SCH2MODEREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH2MODEREG_F2_G);
inv_8044: a_SCH2MODEREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8045: a_EQ1045 <=  n_9138  XOR n_9145;
or2_8046: n_9138 <=  n_9139  OR n_9142;
and2_8047: n_9139 <=  n_9140  AND n_9141;
inv_8048: n_9140  <= TRANSPORT NOT a_N2569_aNOT  ;
delay_8049: n_9141  <= TRANSPORT dbin(4)  ;
and2_8050: n_9142 <=  n_9143  AND n_9144;
delay_8051: n_9143  <= TRANSPORT a_N2569_aNOT  ;
delay_8052: n_9144  <= TRANSPORT a_SCH2MODEREG_F2_G  ;
and1_8053: n_9145 <=  gnd;
delay_8054: n_9146  <= TRANSPORT clk  ;
filter_8055: FILTER_a8237

    PORT MAP (IN1 => n_9146, Y => a_SCH2MODEREG_F2_G_aCLK);
dff_8056: DFF_a8237

    PORT MAP ( D => a_EQ1075, CLK => a_SCH3BAROUT_F0_G_aCLK, CLRN => a_SCH3BAROUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F0_G);
inv_8057: a_SCH3BAROUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8058: a_EQ1075 <=  n_9155  XOR n_9162;
or2_8059: n_9155 <=  n_9156  OR n_9159;
and2_8060: n_9156 <=  n_9157  AND n_9158;
delay_8061: n_9157  <= TRANSPORT a_N2580_aNOT  ;
delay_8062: n_9158  <= TRANSPORT a_SCH3BAROUT_F0_G  ;
and2_8063: n_9159 <=  n_9160  AND n_9161;
inv_8064: n_9160  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_8065: n_9161  <= TRANSPORT dbin(0)  ;
and1_8066: n_9162 <=  gnd;
delay_8067: n_9163  <= TRANSPORT clk  ;
filter_8068: FILTER_a8237

    PORT MAP (IN1 => n_9163, Y => a_SCH3BAROUT_F0_G_aCLK);
dff_8069: DFF_a8237

    PORT MAP ( D => a_EQ1109, CLK => a_SCH3MODEREG_F2_G_aCLK, CLRN => a_SCH3MODEREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH3MODEREG_F2_G);
inv_8070: a_SCH3MODEREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8071: a_EQ1109 <=  n_9171  XOR n_9178;
or2_8072: n_9171 <=  n_9172  OR n_9175;
and2_8073: n_9172 <=  n_9173  AND n_9174;
inv_8074: n_9173  <= TRANSPORT NOT a_N2570_aNOT  ;
delay_8075: n_9174  <= TRANSPORT dbin(4)  ;
and2_8076: n_9175 <=  n_9176  AND n_9177;
delay_8077: n_9176  <= TRANSPORT a_N2570_aNOT  ;
delay_8078: n_9177  <= TRANSPORT a_SCH3MODEREG_F2_G  ;
and1_8079: n_9178 <=  gnd;
delay_8080: n_9179  <= TRANSPORT clk  ;
filter_8081: FILTER_a8237

    PORT MAP (IN1 => n_9179, Y => a_SCH3MODEREG_F2_G_aCLK);
dff_8082: DFF_a8237

    PORT MAP ( D => a_EQ883, CLK => a_SCH0BAROUT_F0_G_aCLK, CLRN => a_SCH0BAROUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F0_G);
inv_8083: a_SCH0BAROUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8084: a_EQ883 <=  n_9188  XOR n_9195;
or2_8085: n_9188 <=  n_9189  OR n_9192;
and2_8086: n_9189 <=  n_9190  AND n_9191;
inv_8087: n_9190  <= TRANSPORT NOT a_N2586  ;
delay_8088: n_9191  <= TRANSPORT a_SCH0BAROUT_F0_G  ;
and2_8089: n_9192 <=  n_9193  AND n_9194;
delay_8090: n_9193  <= TRANSPORT a_N2586  ;
delay_8091: n_9194  <= TRANSPORT dbin(0)  ;
and1_8092: n_9195 <=  gnd;
delay_8093: n_9196  <= TRANSPORT clk  ;
filter_8094: FILTER_a8237

    PORT MAP (IN1 => n_9196, Y => a_SCH0BAROUT_F0_G_aCLK);
delay_8095: a_N2584_aNOT  <= TRANSPORT a_EQ637  ;
xor2_8096: a_EQ637 <=  n_9200  XOR n_9205;
or2_8097: n_9200 <=  n_9201  OR n_9203;
and1_8098: n_9201 <=  n_9202;
delay_8099: n_9202  <= TRANSPORT a_N2352  ;
and1_8100: n_9203 <=  n_9204;
delay_8101: n_9204  <= TRANSPORT a_LC6_D6  ;
and1_8102: n_9205 <=  gnd;
dff_8103: DFF_a8237

    PORT MAP ( D => a_EQ947, CLK => a_SCH1BAROUT_F0_G_aCLK, CLRN => a_SCH1BAROUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F0_G);
inv_8104: a_SCH1BAROUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8105: a_EQ947 <=  n_9213  XOR n_9220;
or2_8106: n_9213 <=  n_9214  OR n_9217;
and2_8107: n_9214 <=  n_9215  AND n_9216;
delay_8108: n_9215  <= TRANSPORT a_N2584_aNOT  ;
delay_8109: n_9216  <= TRANSPORT a_SCH1BAROUT_F0_G  ;
and2_8110: n_9217 <=  n_9218  AND n_9219;
delay_8111: n_9218  <= TRANSPORT dbin(0)  ;
inv_8112: n_9219  <= TRANSPORT NOT a_N2584_aNOT  ;
and1_8113: n_9220 <=  gnd;
delay_8114: n_9221  <= TRANSPORT clk  ;
filter_8115: FILTER_a8237

    PORT MAP (IN1 => n_9221, Y => a_SCH1BAROUT_F0_G_aCLK);
dff_8116: DFF_a8237

    PORT MAP ( D => a_EQ1124, CLK => a_SCOMMANDREG_F1_G_aCLK, CLRN => a_SCOMMANDREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F1_G);
inv_8117: a_SCOMMANDREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8118: a_EQ1124 <=  n_9229  XOR n_9237;
or2_8119: n_9229 <=  n_9230  OR n_9234;
and3_8120: n_9230 <=  n_9231  AND n_9232  AND n_9233;
delay_8121: n_9231  <= TRANSPORT a_N2563_aNOT  ;
delay_8122: n_9232  <= TRANSPORT a_N2571_aNOT  ;
delay_8123: n_9233  <= TRANSPORT a_SCOMMANDREG_F1_G  ;
and2_8124: n_9234 <=  n_9235  AND n_9236;
delay_8125: n_9235  <= TRANSPORT dbin(1)  ;
inv_8126: n_9236  <= TRANSPORT NOT a_N2571_aNOT  ;
and1_8127: n_9237 <=  gnd;
delay_8128: n_9238  <= TRANSPORT clk  ;
filter_8129: FILTER_a8237

    PORT MAP (IN1 => n_9238, Y => a_SCOMMANDREG_F1_G_aCLK);
dff_8130: DFF_a8237

    PORT MAP ( D => a_EQ948, CLK => a_SCH1BAROUT_F1_G_aCLK, CLRN => a_SCH1BAROUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F1_G);
inv_8131: a_SCH1BAROUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8132: a_EQ948 <=  n_9247  XOR n_9254;
or2_8133: n_9247 <=  n_9248  OR n_9251;
and2_8134: n_9248 <=  n_9249  AND n_9250;
delay_8135: n_9249  <= TRANSPORT dbin(1)  ;
inv_8136: n_9250  <= TRANSPORT NOT a_N2584_aNOT  ;
and2_8137: n_9251 <=  n_9252  AND n_9253;
delay_8138: n_9252  <= TRANSPORT a_N2584_aNOT  ;
delay_8139: n_9253  <= TRANSPORT a_SCH1BAROUT_F1_G  ;
and1_8140: n_9254 <=  gnd;
delay_8141: n_9255  <= TRANSPORT clk  ;
filter_8142: FILTER_a8237

    PORT MAP (IN1 => n_9255, Y => a_SCH1BAROUT_F1_G_aCLK);
dff_8143: DFF_a8237

    PORT MAP ( D => a_EQ884, CLK => a_SCH0BAROUT_F1_G_aCLK, CLRN => a_SCH0BAROUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F1_G);
inv_8144: a_SCH0BAROUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8145: a_EQ884 <=  n_9264  XOR n_9271;
or2_8146: n_9264 <=  n_9265  OR n_9268;
and2_8147: n_9265 <=  n_9266  AND n_9267;
delay_8148: n_9266  <= TRANSPORT a_N2586  ;
delay_8149: n_9267  <= TRANSPORT dbin(1)  ;
and2_8150: n_9268 <=  n_9269  AND n_9270;
inv_8151: n_9269  <= TRANSPORT NOT a_N2586  ;
delay_8152: n_9270  <= TRANSPORT a_SCH0BAROUT_F1_G  ;
and1_8153: n_9271 <=  gnd;
delay_8154: n_9272  <= TRANSPORT clk  ;
filter_8155: FILTER_a8237

    PORT MAP (IN1 => n_9272, Y => a_SCH0BAROUT_F1_G_aCLK);
dff_8156: DFF_a8237

    PORT MAP ( D => a_EQ1076, CLK => a_SCH3BAROUT_F1_G_aCLK, CLRN => a_SCH3BAROUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F1_G);
inv_8157: a_SCH3BAROUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8158: a_EQ1076 <=  n_9281  XOR n_9288;
or2_8159: n_9281 <=  n_9282  OR n_9285;
and2_8160: n_9282 <=  n_9283  AND n_9284;
inv_8161: n_9283  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_8162: n_9284  <= TRANSPORT dbin(1)  ;
and2_8163: n_9285 <=  n_9286  AND n_9287;
delay_8164: n_9286  <= TRANSPORT a_N2580_aNOT  ;
delay_8165: n_9287  <= TRANSPORT a_SCH3BAROUT_F1_G  ;
and1_8166: n_9288 <=  gnd;
delay_8167: n_9289  <= TRANSPORT clk  ;
filter_8168: FILTER_a8237

    PORT MAP (IN1 => n_9289, Y => a_SCH3BAROUT_F1_G_aCLK);
dff_8169: DFF_a8237

    PORT MAP ( D => a_EQ949, CLK => a_SCH1BAROUT_F2_G_aCLK, CLRN => a_SCH1BAROUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F2_G);
inv_8170: a_SCH1BAROUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8171: a_EQ949 <=  n_9298  XOR n_9305;
or2_8172: n_9298 <=  n_9299  OR n_9302;
and2_8173: n_9299 <=  n_9300  AND n_9301;
delay_8174: n_9300  <= TRANSPORT dbin(2)  ;
inv_8175: n_9301  <= TRANSPORT NOT a_N2584_aNOT  ;
and2_8176: n_9302 <=  n_9303  AND n_9304;
delay_8177: n_9303  <= TRANSPORT a_N2584_aNOT  ;
delay_8178: n_9304  <= TRANSPORT a_SCH1BAROUT_F2_G  ;
and1_8179: n_9305 <=  gnd;
delay_8180: n_9306  <= TRANSPORT clk  ;
filter_8181: FILTER_a8237

    PORT MAP (IN1 => n_9306, Y => a_SCH1BAROUT_F2_G_aCLK);
dff_8182: DFF_a8237

    PORT MAP ( D => a_EQ1077, CLK => a_SCH3BAROUT_F2_G_aCLK, CLRN => a_SCH3BAROUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F2_G);
inv_8183: a_SCH3BAROUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8184: a_EQ1077 <=  n_9315  XOR n_9322;
or2_8185: n_9315 <=  n_9316  OR n_9319;
and2_8186: n_9316 <=  n_9317  AND n_9318;
inv_8187: n_9317  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_8188: n_9318  <= TRANSPORT dbin(2)  ;
and2_8189: n_9319 <=  n_9320  AND n_9321;
delay_8190: n_9320  <= TRANSPORT a_N2580_aNOT  ;
delay_8191: n_9321  <= TRANSPORT a_SCH3BAROUT_F2_G  ;
and1_8192: n_9322 <=  gnd;
delay_8193: n_9323  <= TRANSPORT clk  ;
filter_8194: FILTER_a8237

    PORT MAP (IN1 => n_9323, Y => a_SCH3BAROUT_F2_G_aCLK);
dff_8195: DFF_a8237

    PORT MAP ( D => a_EQ1013, CLK => a_SCH2BAROUT_F2_G_aCLK, CLRN => a_SCH2BAROUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F2_G);
inv_8196: a_SCH2BAROUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8197: a_EQ1013 <=  n_9332  XOR n_9339;
or2_8198: n_9332 <=  n_9333  OR n_9336;
and2_8199: n_9333 <=  n_9334  AND n_9335;
inv_8200: n_9334  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8201: n_9335  <= TRANSPORT dbin(2)  ;
and2_8202: n_9336 <=  n_9337  AND n_9338;
delay_8203: n_9337  <= TRANSPORT a_N2582_aNOT  ;
delay_8204: n_9338  <= TRANSPORT a_SCH2BAROUT_F2_G  ;
and1_8205: n_9339 <=  gnd;
delay_8206: n_9340  <= TRANSPORT clk  ;
filter_8207: FILTER_a8237

    PORT MAP (IN1 => n_9340, Y => a_SCH2BAROUT_F2_G_aCLK);
dff_8208: DFF_a8237

    PORT MAP ( D => a_EQ885, CLK => a_SCH0BAROUT_F2_G_aCLK, CLRN => a_SCH0BAROUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F2_G);
inv_8209: a_SCH0BAROUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8210: a_EQ885 <=  n_9349  XOR n_9356;
or2_8211: n_9349 <=  n_9350  OR n_9353;
and2_8212: n_9350 <=  n_9351  AND n_9352;
delay_8213: n_9351  <= TRANSPORT a_N2586  ;
delay_8214: n_9352  <= TRANSPORT dbin(2)  ;
and2_8215: n_9353 <=  n_9354  AND n_9355;
inv_8216: n_9354  <= TRANSPORT NOT a_N2586  ;
delay_8217: n_9355  <= TRANSPORT a_SCH0BAROUT_F2_G  ;
and1_8218: n_9356 <=  gnd;
delay_8219: n_9357  <= TRANSPORT clk  ;
filter_8220: FILTER_a8237

    PORT MAP (IN1 => n_9357, Y => a_SCH0BAROUT_F2_G_aCLK);
dff_8221: DFF_a8237

    PORT MAP ( D => a_EQ886, CLK => a_SCH0BAROUT_F3_G_aCLK, CLRN => a_SCH0BAROUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F3_G);
inv_8222: a_SCH0BAROUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8223: a_EQ886 <=  n_9366  XOR n_9373;
or2_8224: n_9366 <=  n_9367  OR n_9370;
and2_8225: n_9367 <=  n_9368  AND n_9369;
delay_8226: n_9368  <= TRANSPORT a_N2586  ;
delay_8227: n_9369  <= TRANSPORT dbin(3)  ;
and2_8228: n_9370 <=  n_9371  AND n_9372;
inv_8229: n_9371  <= TRANSPORT NOT a_N2586  ;
delay_8230: n_9372  <= TRANSPORT a_SCH0BAROUT_F3_G  ;
and1_8231: n_9373 <=  gnd;
delay_8232: n_9374  <= TRANSPORT clk  ;
filter_8233: FILTER_a8237

    PORT MAP (IN1 => n_9374, Y => a_SCH0BAROUT_F3_G_aCLK);
dff_8234: DFF_a8237

    PORT MAP ( D => a_EQ1014, CLK => a_SCH2BAROUT_F3_G_aCLK, CLRN => a_SCH2BAROUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F3_G);
inv_8235: a_SCH2BAROUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8236: a_EQ1014 <=  n_9383  XOR n_9390;
or2_8237: n_9383 <=  n_9384  OR n_9387;
and2_8238: n_9384 <=  n_9385  AND n_9386;
inv_8239: n_9385  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8240: n_9386  <= TRANSPORT dbin(3)  ;
and2_8241: n_9387 <=  n_9388  AND n_9389;
delay_8242: n_9388  <= TRANSPORT a_N2582_aNOT  ;
delay_8243: n_9389  <= TRANSPORT a_SCH2BAROUT_F3_G  ;
and1_8244: n_9390 <=  gnd;
delay_8245: n_9391  <= TRANSPORT clk  ;
filter_8246: FILTER_a8237

    PORT MAP (IN1 => n_9391, Y => a_SCH2BAROUT_F3_G_aCLK);
dff_8247: DFF_a8237

    PORT MAP ( D => a_EQ950, CLK => a_SCH1BAROUT_F3_G_aCLK, CLRN => a_SCH1BAROUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F3_G);
inv_8248: a_SCH1BAROUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8249: a_EQ950 <=  n_9400  XOR n_9407;
or2_8250: n_9400 <=  n_9401  OR n_9404;
and2_8251: n_9401 <=  n_9402  AND n_9403;
delay_8252: n_9402  <= TRANSPORT dbin(3)  ;
inv_8253: n_9403  <= TRANSPORT NOT a_N2584_aNOT  ;
and2_8254: n_9404 <=  n_9405  AND n_9406;
delay_8255: n_9405  <= TRANSPORT a_N2584_aNOT  ;
delay_8256: n_9406  <= TRANSPORT a_SCH1BAROUT_F3_G  ;
and1_8257: n_9407 <=  gnd;
delay_8258: n_9408  <= TRANSPORT clk  ;
filter_8259: FILTER_a8237

    PORT MAP (IN1 => n_9408, Y => a_SCH1BAROUT_F3_G_aCLK);
dff_8260: DFF_a8237

    PORT MAP ( D => a_EQ1078, CLK => a_SCH3BAROUT_F3_G_aCLK, CLRN => a_SCH3BAROUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F3_G);
inv_8261: a_SCH3BAROUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8262: a_EQ1078 <=  n_9417  XOR n_9424;
or2_8263: n_9417 <=  n_9418  OR n_9421;
and2_8264: n_9418 <=  n_9419  AND n_9420;
inv_8265: n_9419  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_8266: n_9420  <= TRANSPORT dbin(3)  ;
and2_8267: n_9421 <=  n_9422  AND n_9423;
delay_8268: n_9422  <= TRANSPORT a_N2580_aNOT  ;
delay_8269: n_9423  <= TRANSPORT a_SCH3BAROUT_F3_G  ;
and1_8270: n_9424 <=  gnd;
delay_8271: n_9425  <= TRANSPORT clk  ;
filter_8272: FILTER_a8237

    PORT MAP (IN1 => n_9425, Y => a_SCH3BAROUT_F3_G_aCLK);
dff_8273: DFF_a8237

    PORT MAP ( D => a_EQ951, CLK => a_SCH1BAROUT_F4_G_aCLK, CLRN => a_SCH1BAROUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F4_G);
inv_8274: a_SCH1BAROUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8275: a_EQ951 <=  n_9434  XOR n_9441;
or2_8276: n_9434 <=  n_9435  OR n_9438;
and2_8277: n_9435 <=  n_9436  AND n_9437;
inv_8278: n_9436  <= TRANSPORT NOT a_N2584_aNOT  ;
delay_8279: n_9437  <= TRANSPORT dbin(4)  ;
and2_8280: n_9438 <=  n_9439  AND n_9440;
delay_8281: n_9439  <= TRANSPORT a_N2584_aNOT  ;
delay_8282: n_9440  <= TRANSPORT a_SCH1BAROUT_F4_G  ;
and1_8283: n_9441 <=  gnd;
delay_8284: n_9442  <= TRANSPORT clk  ;
filter_8285: FILTER_a8237

    PORT MAP (IN1 => n_9442, Y => a_SCH1BAROUT_F4_G_aCLK);
dff_8286: DFF_a8237

    PORT MAP ( D => a_EQ1015, CLK => a_SCH2BAROUT_F4_G_aCLK, CLRN => a_SCH2BAROUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F4_G);
inv_8287: a_SCH2BAROUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8288: a_EQ1015 <=  n_9451  XOR n_9458;
or2_8289: n_9451 <=  n_9452  OR n_9455;
and2_8290: n_9452 <=  n_9453  AND n_9454;
inv_8291: n_9453  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8292: n_9454  <= TRANSPORT dbin(4)  ;
and2_8293: n_9455 <=  n_9456  AND n_9457;
delay_8294: n_9456  <= TRANSPORT a_N2582_aNOT  ;
delay_8295: n_9457  <= TRANSPORT a_SCH2BAROUT_F4_G  ;
and1_8296: n_9458 <=  gnd;
delay_8297: n_9459  <= TRANSPORT clk  ;
filter_8298: FILTER_a8237

    PORT MAP (IN1 => n_9459, Y => a_SCH2BAROUT_F4_G_aCLK);
dff_8299: DFF_a8237

    PORT MAP ( D => a_EQ1079, CLK => a_SCH3BAROUT_F4_G_aCLK, CLRN => a_SCH3BAROUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F4_G);
inv_8300: a_SCH3BAROUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8301: a_EQ1079 <=  n_9468  XOR n_9475;
or2_8302: n_9468 <=  n_9469  OR n_9472;
and2_8303: n_9469 <=  n_9470  AND n_9471;
inv_8304: n_9470  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_8305: n_9471  <= TRANSPORT dbin(4)  ;
and2_8306: n_9472 <=  n_9473  AND n_9474;
delay_8307: n_9473  <= TRANSPORT a_N2580_aNOT  ;
delay_8308: n_9474  <= TRANSPORT a_SCH3BAROUT_F4_G  ;
and1_8309: n_9475 <=  gnd;
delay_8310: n_9476  <= TRANSPORT clk  ;
filter_8311: FILTER_a8237

    PORT MAP (IN1 => n_9476, Y => a_SCH3BAROUT_F4_G_aCLK);
dff_8312: DFF_a8237

    PORT MAP ( D => a_EQ887, CLK => a_SCH0BAROUT_F4_G_aCLK, CLRN => a_SCH0BAROUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F4_G);
inv_8313: a_SCH0BAROUT_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8314: a_EQ887 <=  n_9485  XOR n_9492;
or2_8315: n_9485 <=  n_9486  OR n_9489;
and2_8316: n_9486 <=  n_9487  AND n_9488;
delay_8317: n_9487  <= TRANSPORT a_N2586  ;
delay_8318: n_9488  <= TRANSPORT dbin(4)  ;
and2_8319: n_9489 <=  n_9490  AND n_9491;
inv_8320: n_9490  <= TRANSPORT NOT a_N2586  ;
delay_8321: n_9491  <= TRANSPORT a_SCH0BAROUT_F4_G  ;
and1_8322: n_9492 <=  gnd;
delay_8323: n_9493  <= TRANSPORT clk  ;
filter_8324: FILTER_a8237

    PORT MAP (IN1 => n_9493, Y => a_SCH0BAROUT_F4_G_aCLK);
dff_8325: DFF_a8237

    PORT MAP ( D => a_EQ952, CLK => a_SCH1BAROUT_F5_G_aCLK, CLRN => a_SCH1BAROUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F5_G);
inv_8326: a_SCH1BAROUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8327: a_EQ952 <=  n_9502  XOR n_9509;
or2_8328: n_9502 <=  n_9503  OR n_9506;
and2_8329: n_9503 <=  n_9504  AND n_9505;
inv_8330: n_9504  <= TRANSPORT NOT a_N2584_aNOT  ;
delay_8331: n_9505  <= TRANSPORT dbin(5)  ;
and2_8332: n_9506 <=  n_9507  AND n_9508;
delay_8333: n_9507  <= TRANSPORT a_N2584_aNOT  ;
delay_8334: n_9508  <= TRANSPORT a_SCH1BAROUT_F5_G  ;
and1_8335: n_9509 <=  gnd;
delay_8336: n_9510  <= TRANSPORT clk  ;
filter_8337: FILTER_a8237

    PORT MAP (IN1 => n_9510, Y => a_SCH1BAROUT_F5_G_aCLK);
dff_8338: DFF_a8237

    PORT MAP ( D => a_EQ1016, CLK => a_SCH2BAROUT_F5_G_aCLK, CLRN => a_SCH2BAROUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F5_G);
inv_8339: a_SCH2BAROUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8340: a_EQ1016 <=  n_9519  XOR n_9526;
or2_8341: n_9519 <=  n_9520  OR n_9523;
and2_8342: n_9520 <=  n_9521  AND n_9522;
inv_8343: n_9521  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8344: n_9522  <= TRANSPORT dbin(5)  ;
and2_8345: n_9523 <=  n_9524  AND n_9525;
delay_8346: n_9524  <= TRANSPORT a_N2582_aNOT  ;
delay_8347: n_9525  <= TRANSPORT a_SCH2BAROUT_F5_G  ;
and1_8348: n_9526 <=  gnd;
delay_8349: n_9527  <= TRANSPORT clk  ;
filter_8350: FILTER_a8237

    PORT MAP (IN1 => n_9527, Y => a_SCH2BAROUT_F5_G_aCLK);
dff_8351: DFF_a8237

    PORT MAP ( D => a_EQ888, CLK => a_SCH0BAROUT_F5_G_aCLK, CLRN => a_SCH0BAROUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F5_G);
inv_8352: a_SCH0BAROUT_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8353: a_EQ888 <=  n_9536  XOR n_9543;
or2_8354: n_9536 <=  n_9537  OR n_9540;
and2_8355: n_9537 <=  n_9538  AND n_9539;
delay_8356: n_9538  <= TRANSPORT a_N2586  ;
delay_8357: n_9539  <= TRANSPORT dbin(5)  ;
and2_8358: n_9540 <=  n_9541  AND n_9542;
inv_8359: n_9541  <= TRANSPORT NOT a_N2586  ;
delay_8360: n_9542  <= TRANSPORT a_SCH0BAROUT_F5_G  ;
and1_8361: n_9543 <=  gnd;
delay_8362: n_9544  <= TRANSPORT clk  ;
filter_8363: FILTER_a8237

    PORT MAP (IN1 => n_9544, Y => a_SCH0BAROUT_F5_G_aCLK);
dff_8364: DFF_a8237

    PORT MAP ( D => a_EQ1017, CLK => a_SCH2BAROUT_F6_G_aCLK, CLRN => a_SCH2BAROUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F6_G);
inv_8365: a_SCH2BAROUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8366: a_EQ1017 <=  n_9553  XOR n_9560;
or2_8367: n_9553 <=  n_9554  OR n_9557;
and2_8368: n_9554 <=  n_9555  AND n_9556;
inv_8369: n_9555  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8370: n_9556  <= TRANSPORT dbin(6)  ;
and2_8371: n_9557 <=  n_9558  AND n_9559;
delay_8372: n_9558  <= TRANSPORT a_N2582_aNOT  ;
delay_8373: n_9559  <= TRANSPORT a_SCH2BAROUT_F6_G  ;
and1_8374: n_9560 <=  gnd;
delay_8375: n_9561  <= TRANSPORT clk  ;
filter_8376: FILTER_a8237

    PORT MAP (IN1 => n_9561, Y => a_SCH2BAROUT_F6_G_aCLK);
dff_8377: DFF_a8237

    PORT MAP ( D => a_EQ889, CLK => a_SCH0BAROUT_F6_G_aCLK, CLRN => a_SCH0BAROUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F6_G);
inv_8378: a_SCH0BAROUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8379: a_EQ889 <=  n_9570  XOR n_9577;
or2_8380: n_9570 <=  n_9571  OR n_9574;
and2_8381: n_9571 <=  n_9572  AND n_9573;
delay_8382: n_9572  <= TRANSPORT a_N2586  ;
delay_8383: n_9573  <= TRANSPORT dbin(6)  ;
and2_8384: n_9574 <=  n_9575  AND n_9576;
inv_8385: n_9575  <= TRANSPORT NOT a_N2586  ;
delay_8386: n_9576  <= TRANSPORT a_SCH0BAROUT_F6_G  ;
and1_8387: n_9577 <=  gnd;
delay_8388: n_9578  <= TRANSPORT clk  ;
filter_8389: FILTER_a8237

    PORT MAP (IN1 => n_9578, Y => a_SCH0BAROUT_F6_G_aCLK);
dff_8390: DFF_a8237

    PORT MAP ( D => a_EQ953, CLK => a_SCH1BAROUT_F6_G_aCLK, CLRN => a_SCH1BAROUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F6_G);
inv_8391: a_SCH1BAROUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8392: a_EQ953 <=  n_9587  XOR n_9594;
or2_8393: n_9587 <=  n_9588  OR n_9591;
and2_8394: n_9588 <=  n_9589  AND n_9590;
delay_8395: n_9589  <= TRANSPORT dbin(6)  ;
inv_8396: n_9590  <= TRANSPORT NOT a_N2584_aNOT  ;
and2_8397: n_9591 <=  n_9592  AND n_9593;
delay_8398: n_9592  <= TRANSPORT a_N2584_aNOT  ;
delay_8399: n_9593  <= TRANSPORT a_SCH1BAROUT_F6_G  ;
and1_8400: n_9594 <=  gnd;
delay_8401: n_9595  <= TRANSPORT clk  ;
filter_8402: FILTER_a8237

    PORT MAP (IN1 => n_9595, Y => a_SCH1BAROUT_F6_G_aCLK);
dff_8403: DFF_a8237

    PORT MAP ( D => a_EQ1081, CLK => a_SCH3BAROUT_F6_G_aCLK, CLRN => a_SCH3BAROUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH3BAROUT_F6_G);
inv_8404: a_SCH3BAROUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8405: a_EQ1081 <=  n_9604  XOR n_9611;
or2_8406: n_9604 <=  n_9605  OR n_9608;
and2_8407: n_9605 <=  n_9606  AND n_9607;
inv_8408: n_9606  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_8409: n_9607  <= TRANSPORT dbin(6)  ;
and2_8410: n_9608 <=  n_9609  AND n_9610;
delay_8411: n_9609  <= TRANSPORT a_N2580_aNOT  ;
delay_8412: n_9610  <= TRANSPORT a_SCH3BAROUT_F6_G  ;
and1_8413: n_9611 <=  gnd;
delay_8414: n_9612  <= TRANSPORT clk  ;
filter_8415: FILTER_a8237

    PORT MAP (IN1 => n_9612, Y => a_SCH3BAROUT_F6_G_aCLK);
dff_8416: DFF_a8237

    PORT MAP ( D => a_EQ1018, CLK => a_SCH2BAROUT_F7_G_aCLK, CLRN => a_SCH2BAROUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH2BAROUT_F7_G);
inv_8417: a_SCH2BAROUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8418: a_EQ1018 <=  n_9621  XOR n_9628;
or2_8419: n_9621 <=  n_9622  OR n_9625;
and2_8420: n_9622 <=  n_9623  AND n_9624;
inv_8421: n_9623  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_8422: n_9624  <= TRANSPORT dbin(7)  ;
and2_8423: n_9625 <=  n_9626  AND n_9627;
delay_8424: n_9626  <= TRANSPORT a_N2582_aNOT  ;
delay_8425: n_9627  <= TRANSPORT a_SCH2BAROUT_F7_G  ;
and1_8426: n_9628 <=  gnd;
delay_8427: n_9629  <= TRANSPORT clk  ;
filter_8428: FILTER_a8237

    PORT MAP (IN1 => n_9629, Y => a_SCH2BAROUT_F7_G_aCLK);
dff_8429: DFF_a8237

    PORT MAP ( D => a_EQ917, CLK => a_SCH0MODEREG_F2_G_aCLK, CLRN => a_SCH0MODEREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH0MODEREG_F2_G);
inv_8430: a_SCH0MODEREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8431: a_EQ917 <=  n_9637  XOR n_9644;
or2_8432: n_9637 <=  n_9638  OR n_9641;
and2_8433: n_9638 <=  n_9639  AND n_9640;
inv_8434: n_9639  <= TRANSPORT NOT a_N2567  ;
delay_8435: n_9640  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and2_8436: n_9641 <=  n_9642  AND n_9643;
delay_8437: n_9642  <= TRANSPORT a_N2567  ;
delay_8438: n_9643  <= TRANSPORT dbin(4)  ;
and1_8439: n_9644 <=  gnd;
delay_8440: n_9645  <= TRANSPORT clk  ;
filter_8441: FILTER_a8237

    PORT MAP (IN1 => n_9645, Y => a_SCH0MODEREG_F2_G_aCLK);
dff_8442: DFF_a8237

    PORT MAP ( D => a_EQ890, CLK => a_SCH0BAROUT_F7_G_aCLK, CLRN => a_SCH0BAROUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH0BAROUT_F7_G);
inv_8443: a_SCH0BAROUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8444: a_EQ890 <=  n_9654  XOR n_9661;
or2_8445: n_9654 <=  n_9655  OR n_9658;
and2_8446: n_9655 <=  n_9656  AND n_9657;
delay_8447: n_9656  <= TRANSPORT a_N2586  ;
delay_8448: n_9657  <= TRANSPORT dbin(7)  ;
and2_8449: n_9658 <=  n_9659  AND n_9660;
inv_8450: n_9659  <= TRANSPORT NOT a_N2586  ;
delay_8451: n_9660  <= TRANSPORT a_SCH0BAROUT_F7_G  ;
and1_8452: n_9661 <=  gnd;
delay_8453: n_9662  <= TRANSPORT clk  ;
filter_8454: FILTER_a8237

    PORT MAP (IN1 => n_9662, Y => a_SCH0BAROUT_F7_G_aCLK);
dff_8455: DFF_a8237

    PORT MAP ( D => a_EQ981, CLK => a_SCH1MODEREG_F2_G_aCLK, CLRN => a_SCH1MODEREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH1MODEREG_F2_G);
inv_8456: a_SCH1MODEREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8457: a_EQ981 <=  n_9670  XOR n_9677;
or2_8458: n_9670 <=  n_9671  OR n_9674;
and2_8459: n_9671 <=  n_9672  AND n_9673;
inv_8460: n_9672  <= TRANSPORT NOT a_N2568  ;
delay_8461: n_9673  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and2_8462: n_9674 <=  n_9675  AND n_9676;
delay_8463: n_9675  <= TRANSPORT a_N2568  ;
delay_8464: n_9676  <= TRANSPORT dbin(4)  ;
and1_8465: n_9677 <=  gnd;
delay_8466: n_9678  <= TRANSPORT clk  ;
filter_8467: FILTER_a8237

    PORT MAP (IN1 => n_9678, Y => a_SCH1MODEREG_F2_G_aCLK);
dff_8468: DFF_a8237

    PORT MAP ( D => a_EQ954, CLK => a_SCH1BAROUT_F7_G_aCLK, CLRN => a_SCH1BAROUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH1BAROUT_F7_G);
inv_8469: a_SCH1BAROUT_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8470: a_EQ954 <=  n_9687  XOR n_9694;
or2_8471: n_9687 <=  n_9688  OR n_9691;
and2_8472: n_9688 <=  n_9689  AND n_9690;
inv_8473: n_9689  <= TRANSPORT NOT a_N2584_aNOT  ;
delay_8474: n_9690  <= TRANSPORT dbin(7)  ;
and2_8475: n_9691 <=  n_9692  AND n_9693;
delay_8476: n_9692  <= TRANSPORT a_N2584_aNOT  ;
delay_8477: n_9693  <= TRANSPORT a_SCH1BAROUT_F7_G  ;
and1_8478: n_9694 <=  gnd;
delay_8479: n_9695  <= TRANSPORT clk  ;
filter_8480: FILTER_a8237

    PORT MAP (IN1 => n_9695, Y => a_SCH1BAROUT_F7_G_aCLK);
dff_8481: DFF_a8237

    PORT MAP ( D => a_EQ1043, CLK => a_SCH2MODEREG_F0_G_aCLK, CLRN => a_SCH2MODEREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH2MODEREG_F0_G);
inv_8482: a_SCH2MODEREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8483: a_EQ1043 <=  n_9703  XOR n_9710;
or2_8484: n_9703 <=  n_9704  OR n_9707;
and2_8485: n_9704 <=  n_9705  AND n_9706;
delay_8486: n_9705  <= TRANSPORT a_N2569_aNOT  ;
delay_8487: n_9706  <= TRANSPORT a_SCH2MODEREG_F0_G  ;
and2_8488: n_9707 <=  n_9708  AND n_9709;
inv_8489: n_9708  <= TRANSPORT NOT a_N2569_aNOT  ;
delay_8490: n_9709  <= TRANSPORT dbin(2)  ;
and1_8491: n_9710 <=  gnd;
delay_8492: n_9711  <= TRANSPORT clk  ;
filter_8493: FILTER_a8237

    PORT MAP (IN1 => n_9711, Y => a_SCH2MODEREG_F0_G_aCLK);
dff_8494: DFF_a8237

    PORT MAP ( D => a_EQ979, CLK => a_SCH1MODEREG_F0_G_aCLK, CLRN => a_SCH1MODEREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH1MODEREG_F0_G);
inv_8495: a_SCH1MODEREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8496: a_EQ979 <=  n_9719  XOR n_9726;
or2_8497: n_9719 <=  n_9720  OR n_9723;
and2_8498: n_9720 <=  n_9721  AND n_9722;
inv_8499: n_9721  <= TRANSPORT NOT a_N2568  ;
delay_8500: n_9722  <= TRANSPORT a_SCH1MODEREG_F0_G  ;
and2_8501: n_9723 <=  n_9724  AND n_9725;
delay_8502: n_9724  <= TRANSPORT a_N2568  ;
delay_8503: n_9725  <= TRANSPORT dbin(2)  ;
and1_8504: n_9726 <=  gnd;
delay_8505: n_9727  <= TRANSPORT clk  ;
filter_8506: FILTER_a8237

    PORT MAP (IN1 => n_9727, Y => a_SCH1MODEREG_F0_G_aCLK);
dff_8507: DFF_a8237

    PORT MAP ( D => a_EQ915, CLK => a_SCH0MODEREG_F0_G_aCLK, CLRN => a_SCH0MODEREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH0MODEREG_F0_G);
inv_8508: a_SCH0MODEREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8509: a_EQ915 <=  n_9735  XOR n_9742;
or2_8510: n_9735 <=  n_9736  OR n_9739;
and2_8511: n_9736 <=  n_9737  AND n_9738;
inv_8512: n_9737  <= TRANSPORT NOT a_N2567  ;
delay_8513: n_9738  <= TRANSPORT a_SCH0MODEREG_F0_G  ;
and2_8514: n_9739 <=  n_9740  AND n_9741;
delay_8515: n_9740  <= TRANSPORT a_N2567  ;
delay_8516: n_9741  <= TRANSPORT dbin(2)  ;
and1_8517: n_9742 <=  gnd;
delay_8518: n_9743  <= TRANSPORT clk  ;
filter_8519: FILTER_a8237

    PORT MAP (IN1 => n_9743, Y => a_SCH0MODEREG_F0_G_aCLK);
dff_8520: DFF_a8237

    PORT MAP ( D => a_EQ1107, CLK => a_SCH3MODEREG_F0_G_aCLK, CLRN => a_SCH3MODEREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH3MODEREG_F0_G);
inv_8521: a_SCH3MODEREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8522: a_EQ1107 <=  n_9751  XOR n_9758;
or2_8523: n_9751 <=  n_9752  OR n_9755;
and2_8524: n_9752 <=  n_9753  AND n_9754;
delay_8525: n_9753  <= TRANSPORT a_N2570_aNOT  ;
delay_8526: n_9754  <= TRANSPORT a_SCH3MODEREG_F0_G  ;
and2_8527: n_9755 <=  n_9756  AND n_9757;
inv_8528: n_9756  <= TRANSPORT NOT a_N2570_aNOT  ;
delay_8529: n_9757  <= TRANSPORT dbin(2)  ;
and1_8530: n_9758 <=  gnd;
delay_8531: n_9759  <= TRANSPORT clk  ;
filter_8532: FILTER_a8237

    PORT MAP (IN1 => n_9759, Y => a_SCH3MODEREG_F0_G_aCLK);
dff_8533: DFF_a8237

    PORT MAP ( D => a_EQ980, CLK => a_SCH1MODEREG_F1_G_aCLK, CLRN => a_SCH1MODEREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH1MODEREG_F1_G);
inv_8534: a_SCH1MODEREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8535: a_EQ980 <=  n_9767  XOR n_9774;
or2_8536: n_9767 <=  n_9768  OR n_9771;
and2_8537: n_9768 <=  n_9769  AND n_9770;
inv_8538: n_9769  <= TRANSPORT NOT a_N2568  ;
delay_8539: n_9770  <= TRANSPORT a_SCH1MODEREG_F1_G  ;
and2_8540: n_9771 <=  n_9772  AND n_9773;
delay_8541: n_9772  <= TRANSPORT a_N2568  ;
delay_8542: n_9773  <= TRANSPORT dbin(3)  ;
and1_8543: n_9774 <=  gnd;
delay_8544: n_9775  <= TRANSPORT clk  ;
filter_8545: FILTER_a8237

    PORT MAP (IN1 => n_9775, Y => a_SCH1MODEREG_F1_G_aCLK);
dff_8546: DFF_a8237

    PORT MAP ( D => a_EQ1108, CLK => a_SCH3MODEREG_F1_G_aCLK, CLRN => a_SCH3MODEREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH3MODEREG_F1_G);
inv_8547: a_SCH3MODEREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8548: a_EQ1108 <=  n_9783  XOR n_9790;
or2_8549: n_9783 <=  n_9784  OR n_9787;
and2_8550: n_9784 <=  n_9785  AND n_9786;
delay_8551: n_9785  <= TRANSPORT a_N2570_aNOT  ;
delay_8552: n_9786  <= TRANSPORT a_SCH3MODEREG_F1_G  ;
and2_8553: n_9787 <=  n_9788  AND n_9789;
inv_8554: n_9788  <= TRANSPORT NOT a_N2570_aNOT  ;
delay_8555: n_9789  <= TRANSPORT dbin(3)  ;
and1_8556: n_9790 <=  gnd;
delay_8557: n_9791  <= TRANSPORT clk  ;
filter_8558: FILTER_a8237

    PORT MAP (IN1 => n_9791, Y => a_SCH3MODEREG_F1_G_aCLK);
dff_8559: DFF_a8237

    PORT MAP ( D => a_EQ916, CLK => a_SCH0MODEREG_F1_G_aCLK, CLRN => a_SCH0MODEREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH0MODEREG_F1_G);
inv_8560: a_SCH0MODEREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8561: a_EQ916 <=  n_9799  XOR n_9806;
or2_8562: n_9799 <=  n_9800  OR n_9803;
and2_8563: n_9800 <=  n_9801  AND n_9802;
inv_8564: n_9801  <= TRANSPORT NOT a_N2567  ;
delay_8565: n_9802  <= TRANSPORT a_SCH0MODEREG_F1_G  ;
and2_8566: n_9803 <=  n_9804  AND n_9805;
delay_8567: n_9804  <= TRANSPORT a_N2567  ;
delay_8568: n_9805  <= TRANSPORT dbin(3)  ;
and1_8569: n_9806 <=  gnd;
delay_8570: n_9807  <= TRANSPORT clk  ;
filter_8571: FILTER_a8237

    PORT MAP (IN1 => n_9807, Y => a_SCH0MODEREG_F1_G_aCLK);
dff_8572: DFF_a8237

    PORT MAP ( D => a_EQ1044, CLK => a_SCH2MODEREG_F1_G_aCLK, CLRN => a_SCH2MODEREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH2MODEREG_F1_G);
inv_8573: a_SCH2MODEREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8574: a_EQ1044 <=  n_9815  XOR n_9822;
or2_8575: n_9815 <=  n_9816  OR n_9819;
and2_8576: n_9816 <=  n_9817  AND n_9818;
delay_8577: n_9817  <= TRANSPORT a_N2569_aNOT  ;
delay_8578: n_9818  <= TRANSPORT a_SCH2MODEREG_F1_G  ;
and2_8579: n_9819 <=  n_9820  AND n_9821;
inv_8580: n_9820  <= TRANSPORT NOT a_N2569_aNOT  ;
delay_8581: n_9821  <= TRANSPORT dbin(3)  ;
and1_8582: n_9822 <=  gnd;
delay_8583: n_9823  <= TRANSPORT clk  ;
filter_8584: FILTER_a8237

    PORT MAP (IN1 => n_9823, Y => a_SCH2MODEREG_F1_G_aCLK);
delay_8585: a_LC2_E21  <= TRANSPORT a_EQ375  ;
xor2_8586: a_EQ375 <=  n_9827  XOR n_9834;
or2_8587: n_9827 <=  n_9828  OR n_9831;
and2_8588: n_9828 <=  n_9829  AND n_9830;
inv_8589: n_9829  <= TRANSPORT NOT a_N2376  ;
delay_8590: n_9830  <= TRANSPORT a_SH2WRDCNTREG_F10_G  ;
and2_8591: n_9831 <=  n_9832  AND n_9833;
inv_8592: n_9832  <= TRANSPORT NOT a_N2377  ;
delay_8593: n_9833  <= TRANSPORT a_SH3WRDCNTREG_F10_G  ;
and1_8594: n_9834 <=  gnd;
delay_8595: a_N1162_aNOT  <= TRANSPORT a_EQ372  ;
xor2_8596: a_EQ372 <=  n_9837  XOR n_9848;
or3_8597: n_9837 <=  n_9838  OR n_9841  OR n_9844;
and2_8598: n_9838 <=  n_9839  AND n_9840;
inv_8599: n_9839  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
delay_8600: n_9840  <= TRANSPORT a_N3546  ;
and2_8601: n_9841 <=  n_9842  AND n_9843;
inv_8602: n_9842  <= TRANSPORT NOT a_N2557  ;
delay_8603: n_9843  <= TRANSPORT a_N3546  ;
and3_8604: n_9844 <=  n_9845  AND n_9846  AND n_9847;
delay_8605: n_9845  <= TRANSPORT a_N2557  ;
delay_8606: n_9846  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_8607: n_9847  <= TRANSPORT NOT a_N3546  ;
and1_8608: n_9848 <=  gnd;
delay_8609: a_N1168  <= TRANSPORT a_EQ377  ;
xor2_8610: a_EQ377 <=  n_9851  XOR n_9858;
or2_8611: n_9851 <=  n_9852  OR n_9855;
and2_8612: n_9852 <=  n_9853  AND n_9854;
delay_8613: n_9853  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_8614: n_9854  <= TRANSPORT a_SH1WRDCNTREG_F10_G  ;
and2_8615: n_9855 <=  n_9856  AND n_9857;
inv_8616: n_9856  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_8617: n_9857  <= TRANSPORT a_SH0WRDCNTREG_F10_G  ;
and1_8618: n_9858 <=  gnd;
delay_8619: a_N1169  <= TRANSPORT a_EQ378  ;
xor2_8620: a_EQ378 <=  n_9861  XOR n_9870;
or3_8621: n_9861 <=  n_9862  OR n_9864  OR n_9867;
and1_8622: n_9862 <=  n_9863;
delay_8623: n_9863  <= TRANSPORT startdma  ;
and2_8624: n_9864 <=  n_9865  AND n_9866;
inv_8625: n_9865  <= TRANSPORT NOT a_N2531  ;
delay_8626: n_9866  <= TRANSPORT a_N1162_aNOT  ;
and2_8627: n_9867 <=  n_9868  AND n_9869;
delay_8628: n_9868  <= TRANSPORT a_N2531  ;
delay_8629: n_9869  <= TRANSPORT a_N1168  ;
and1_8630: n_9870 <=  gnd;
delay_8631: a_LC3_E21  <= TRANSPORT a_EQ376  ;
xor2_8632: a_EQ376 <=  n_9873  XOR n_9880;
or2_8633: n_9873 <=  n_9874  OR n_9877;
and2_8634: n_9874 <=  n_9875  AND n_9876;
inv_8635: n_9875  <= TRANSPORT NOT a_N88_aNOT  ;
delay_8636: n_9876  <= TRANSPORT a_SH1WRDCNTREG_F10_G  ;
and2_8637: n_9877 <=  n_9878  AND n_9879;
inv_8638: n_9878  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_8639: n_9879  <= TRANSPORT a_SH0WRDCNTREG_F10_G  ;
and1_8640: n_9880 <=  gnd;
dff_8641: DFF_a8237

    PORT MAP ( D => a_EQ842, CLK => a_N3546_aCLK, CLRN => a_N3546_aCLRN, PRN => vcc,
          Q => a_N3546);
inv_8642: a_N3546_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8643: a_EQ842 <=  n_9887  XOR n_9897;
or3_8644: n_9887 <=  n_9888  OR n_9891  OR n_9894;
and2_8645: n_9888 <=  n_9889  AND n_9890;
delay_8646: n_9889  <= TRANSPORT a_LC2_E21  ;
delay_8647: n_9890  <= TRANSPORT a_N1169  ;
and2_8648: n_9891 <=  n_9892  AND n_9893;
delay_8649: n_9892  <= TRANSPORT a_N1169  ;
inv_8650: n_9893  <= TRANSPORT NOT startdma  ;
and2_8651: n_9894 <=  n_9895  AND n_9896;
delay_8652: n_9895  <= TRANSPORT a_N1169  ;
delay_8653: n_9896  <= TRANSPORT a_LC3_E21  ;
and1_8654: n_9897 <=  gnd;
delay_8655: n_9898  <= TRANSPORT clk  ;
filter_8656: FILTER_a8237

    PORT MAP (IN1 => n_9898, Y => a_N3546_aCLK);
delay_8657: a_LC4_A20  <= TRANSPORT a_EQ259  ;
xor2_8658: a_EQ259 <=  n_9902  XOR n_9917;
or4_8659: n_9902 <=  n_9903  OR n_9906  OR n_9909  OR n_9912;
and2_8660: n_9903 <=  n_9904  AND n_9905;
inv_8661: n_9904  <= TRANSPORT NOT a_LC4_A13_aNOT  ;
delay_8662: n_9905  <= TRANSPORT a_N3545  ;
and2_8663: n_9906 <=  n_9907  AND n_9908;
inv_8664: n_9907  <= TRANSPORT NOT a_N2557  ;
delay_8665: n_9908  <= TRANSPORT a_N3545  ;
and2_8666: n_9909 <=  n_9910  AND n_9911;
delay_8667: n_9910  <= TRANSPORT a_N3546  ;
delay_8668: n_9911  <= TRANSPORT a_N3545  ;
and4_8669: n_9912 <=  n_9913  AND n_9914  AND n_9915  AND n_9916;
delay_8670: n_9913  <= TRANSPORT a_N2557  ;
delay_8671: n_9914  <= TRANSPORT a_LC4_A13_aNOT  ;
inv_8672: n_9915  <= TRANSPORT NOT a_N3546  ;
inv_8673: n_9916  <= TRANSPORT NOT a_N3545  ;
and1_8674: n_9917 <=  gnd;
delay_8675: a_LC2_A20  <= TRANSPORT a_EQ258  ;
xor2_8676: a_EQ258 <=  n_9920  XOR n_9927;
or2_8677: n_9920 <=  n_9921  OR n_9924;
and2_8678: n_9921 <=  n_9922  AND n_9923;
delay_8679: n_9922  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_8680: n_9923  <= TRANSPORT a_SH1WRDCNTREG_F11_G  ;
and2_8681: n_9924 <=  n_9925  AND n_9926;
inv_8682: n_9925  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_8683: n_9926  <= TRANSPORT a_SH0WRDCNTREG_F11_G  ;
and1_8684: n_9927 <=  gnd;
delay_8685: a_N517_aNOT  <= TRANSPORT a_EQ262  ;
xor2_8686: a_EQ262 <=  n_9930  XOR n_9937;
or2_8687: n_9930 <=  n_9931  OR n_9934;
and2_8688: n_9931 <=  n_9932  AND n_9933;
inv_8689: n_9932  <= TRANSPORT NOT a_N2531  ;
delay_8690: n_9933  <= TRANSPORT a_LC4_A20  ;
and2_8691: n_9934 <=  n_9935  AND n_9936;
delay_8692: n_9935  <= TRANSPORT a_N2531  ;
delay_8693: n_9936  <= TRANSPORT a_LC2_A20  ;
and1_8694: n_9937 <=  gnd;
delay_8695: a_LC8_A26  <= TRANSPORT a_EQ261  ;
xor2_8696: a_EQ261 <=  n_9940  XOR n_9947;
or2_8697: n_9940 <=  n_9941  OR n_9944;
and2_8698: n_9941 <=  n_9942  AND n_9943;
inv_8699: n_9942  <= TRANSPORT NOT a_N2377  ;
delay_8700: n_9943  <= TRANSPORT a_SH3WRDCNTREG_F11_G  ;
and2_8701: n_9944 <=  n_9945  AND n_9946;
inv_8702: n_9945  <= TRANSPORT NOT a_N88_aNOT  ;
delay_8703: n_9946  <= TRANSPORT a_SH1WRDCNTREG_F11_G  ;
and1_8704: n_9947 <=  gnd;
delay_8705: a_LC8_A20  <= TRANSPORT a_EQ260  ;
xor2_8706: a_EQ260 <=  n_9950  XOR n_9957;
or2_8707: n_9950 <=  n_9951  OR n_9954;
and2_8708: n_9951 <=  n_9952  AND n_9953;
inv_8709: n_9952  <= TRANSPORT NOT a_N2376  ;
delay_8710: n_9953  <= TRANSPORT a_SH2WRDCNTREG_F11_G  ;
and2_8711: n_9954 <=  n_9955  AND n_9956;
inv_8712: n_9955  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_8713: n_9956  <= TRANSPORT a_SH0WRDCNTREG_F11_G  ;
and1_8714: n_9957 <=  gnd;
dff_8715: DFF_a8237

    PORT MAP ( D => a_EQ841, CLK => a_N3545_aCLK, CLRN => a_N3545_aCLRN, PRN => vcc,
          Q => a_N3545);
inv_8716: a_N3545_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8717: a_EQ841 <=  n_9964  XOR n_9974;
or3_8718: n_9964 <=  n_9965  OR n_9968  OR n_9971;
and2_8719: n_9965 <=  n_9966  AND n_9967;
delay_8720: n_9966  <= TRANSPORT a_N517_aNOT  ;
inv_8721: n_9967  <= TRANSPORT NOT startdma  ;
and2_8722: n_9968 <=  n_9969  AND n_9970;
delay_8723: n_9969  <= TRANSPORT a_LC8_A26  ;
delay_8724: n_9970  <= TRANSPORT startdma  ;
and2_8725: n_9971 <=  n_9972  AND n_9973;
delay_8726: n_9972  <= TRANSPORT a_LC8_A20  ;
delay_8727: n_9973  <= TRANSPORT startdma  ;
and1_8728: n_9974 <=  gnd;
delay_8729: n_9975  <= TRANSPORT clk  ;
filter_8730: FILTER_a8237

    PORT MAP (IN1 => n_9975, Y => a_N3545_aCLK);
delay_8731: a_LC3_A1  <= TRANSPORT a_EQ403  ;
xor2_8732: a_EQ403 <=  n_9979  XOR n_9986;
or2_8733: n_9979 <=  n_9980  OR n_9983;
and2_8734: n_9980 <=  n_9981  AND n_9982;
inv_8735: n_9981  <= TRANSPORT NOT a_N2377  ;
delay_8736: n_9982  <= TRANSPORT a_SH3WRDCNTREG_F12_G  ;
and2_8737: n_9983 <=  n_9984  AND n_9985;
inv_8738: n_9984  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_8739: n_9985  <= TRANSPORT a_SH0WRDCNTREG_F12_G  ;
and1_8740: n_9986 <=  gnd;
delay_8741: a_N1297_aNOT  <= TRANSPORT a_EQ410  ;
xor2_8742: a_EQ410 <=  n_9989  XOR n_9996;
or2_8743: n_9989 <=  n_9990  OR n_9993;
and2_8744: n_9990 <=  n_9991  AND n_9992;
delay_8745: n_9991  <= TRANSPORT a_N2557  ;
inv_8746: n_9992  <= TRANSPORT NOT a_LC6_A20  ;
and2_8747: n_9993 <=  n_9994  AND n_9995;
inv_8748: n_9994  <= TRANSPORT NOT a_N2557  ;
delay_8749: n_9995  <= TRANSPORT a_N3544  ;
and1_8750: n_9996 <=  gnd;
delay_8751: a_N1286  <= TRANSPORT a_EQ402  ;
xor2_8752: a_EQ402 <=  n_9999  XOR n_10006;
or2_8753: n_9999 <=  n_10000  OR n_10003;
and2_8754: n_10000 <=  n_10001  AND n_10002;
inv_8755: n_10001  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_8756: n_10002  <= TRANSPORT a_SH0WRDCNTREG_F12_G  ;
and2_8757: n_10003 <=  n_10004  AND n_10005;
delay_8758: n_10004  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_8759: n_10005  <= TRANSPORT a_SH1WRDCNTREG_F12_G  ;
and1_8760: n_10006 <=  gnd;
delay_8761: a_N1285  <= TRANSPORT a_EQ401  ;
xor2_8762: a_EQ401 <=  n_10009  XOR n_10018;
or3_8763: n_10009 <=  n_10010  OR n_10012  OR n_10015;
and1_8764: n_10010 <=  n_10011;
delay_8765: n_10011  <= TRANSPORT startdma  ;
and2_8766: n_10012 <=  n_10013  AND n_10014;
inv_8767: n_10013  <= TRANSPORT NOT a_N2531  ;
delay_8768: n_10014  <= TRANSPORT a_N1297_aNOT  ;
and2_8769: n_10015 <=  n_10016  AND n_10017;
delay_8770: n_10016  <= TRANSPORT a_N2531  ;
delay_8771: n_10017  <= TRANSPORT a_N1286  ;
and1_8772: n_10018 <=  gnd;
delay_8773: a_LC1_A1  <= TRANSPORT a_EQ404  ;
xor2_8774: a_EQ404 <=  n_10021  XOR n_10028;
or2_8775: n_10021 <=  n_10022  OR n_10025;
and2_8776: n_10022 <=  n_10023  AND n_10024;
inv_8777: n_10023  <= TRANSPORT NOT a_N2376  ;
delay_8778: n_10024  <= TRANSPORT a_SH2WRDCNTREG_F12_G  ;
and2_8779: n_10025 <=  n_10026  AND n_10027;
inv_8780: n_10026  <= TRANSPORT NOT a_N88_aNOT  ;
delay_8781: n_10027  <= TRANSPORT a_SH1WRDCNTREG_F12_G  ;
and1_8782: n_10028 <=  gnd;
dff_8783: DFF_a8237

    PORT MAP ( D => a_EQ840, CLK => a_N3544_aCLK, CLRN => a_N3544_aCLRN, PRN => vcc,
          Q => a_N3544);
inv_8784: a_N3544_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8785: a_EQ840 <=  n_10035  XOR n_10045;
or3_8786: n_10035 <=  n_10036  OR n_10039  OR n_10042;
and2_8787: n_10036 <=  n_10037  AND n_10038;
delay_8788: n_10037  <= TRANSPORT a_LC3_A1  ;
delay_8789: n_10038  <= TRANSPORT a_N1285  ;
and2_8790: n_10039 <=  n_10040  AND n_10041;
delay_8791: n_10040  <= TRANSPORT a_N1285  ;
inv_8792: n_10041  <= TRANSPORT NOT startdma  ;
and2_8793: n_10042 <=  n_10043  AND n_10044;
delay_8794: n_10043  <= TRANSPORT a_N1285  ;
delay_8795: n_10044  <= TRANSPORT a_LC1_A1  ;
and1_8796: n_10045 <=  gnd;
delay_8797: n_10046  <= TRANSPORT clk  ;
filter_8798: FILTER_a8237

    PORT MAP (IN1 => n_10046, Y => a_N3544_aCLK);
delay_8799: a_LC7_E14  <= TRANSPORT a_EQ340  ;
xor2_8800: a_EQ340 <=  n_10051  XOR n_10058;
or2_8801: n_10051 <=  n_10052  OR n_10055;
and2_8802: n_10052 <=  n_10053  AND n_10054;
delay_8803: n_10053  <= TRANSPORT a_N2557  ;
delay_8804: n_10054  <= TRANSPORT a_N2594_aNOT  ;
and2_8805: n_10055 <=  n_10056  AND n_10057;
inv_8806: n_10056  <= TRANSPORT NOT a_N2557  ;
delay_8807: n_10057  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and1_8808: n_10058 <=  gnd;
delay_8809: a_LC4_E14  <= TRANSPORT a_EQ339  ;
xor2_8810: a_EQ339 <=  n_10061  XOR n_10068;
or2_8811: n_10061 <=  n_10062  OR n_10065;
and2_8812: n_10062 <=  n_10063  AND n_10064;
delay_8813: n_10063  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_8814: n_10064  <= TRANSPORT a_SCH1ADDRREG_F13_G  ;
and2_8815: n_10065 <=  n_10066  AND n_10067;
inv_8816: n_10066  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_8817: n_10067  <= TRANSPORT a_SCH0ADDRREG_F13_G  ;
and1_8818: n_10068 <=  gnd;
delay_8819: a_N1019_aNOT  <= TRANSPORT a_EQ341  ;
xor2_8820: a_EQ341 <=  n_10071  XOR n_10078;
or2_8821: n_10071 <=  n_10072  OR n_10075;
and2_8822: n_10072 <=  n_10073  AND n_10074;
inv_8823: n_10073  <= TRANSPORT NOT a_N2531  ;
delay_8824: n_10074  <= TRANSPORT a_LC7_E14  ;
and2_8825: n_10075 <=  n_10076  AND n_10077;
delay_8826: n_10076  <= TRANSPORT a_N2531  ;
delay_8827: n_10077  <= TRANSPORT a_LC4_E14  ;
and1_8828: n_10078 <=  gnd;
delay_8829: a_LC5_E14  <= TRANSPORT a_EQ338  ;
xor2_8830: a_EQ338 <=  n_10081  XOR n_10088;
or2_8831: n_10081 <=  n_10082  OR n_10085;
and2_8832: n_10082 <=  n_10083  AND n_10084;
inv_8833: n_10083  <= TRANSPORT NOT a_N2377  ;
delay_8834: n_10084  <= TRANSPORT a_SCH3ADDRREG_F13_G  ;
and2_8835: n_10085 <=  n_10086  AND n_10087;
inv_8836: n_10086  <= TRANSPORT NOT a_N88_aNOT  ;
delay_8837: n_10087  <= TRANSPORT a_SCH1ADDRREG_F13_G  ;
and1_8838: n_10088 <=  gnd;
delay_8839: a_LC6_E14  <= TRANSPORT a_EQ337  ;
xor2_8840: a_EQ337 <=  n_10091  XOR n_10098;
or2_8841: n_10091 <=  n_10092  OR n_10095;
and2_8842: n_10092 <=  n_10093  AND n_10094;
inv_8843: n_10093  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_8844: n_10094  <= TRANSPORT a_SCH0ADDRREG_F13_G  ;
and2_8845: n_10095 <=  n_10096  AND n_10097;
inv_8846: n_10096  <= TRANSPORT NOT a_N2376  ;
delay_8847: n_10097  <= TRANSPORT a_SCH2ADDRREG_F13_G  ;
and1_8848: n_10098 <=  gnd;
dff_8849: DFF_a8237

    PORT MAP ( D => a_EQ859, CLK => a_SADDRESSOUT_F13_G_aCLK, CLRN => a_SADDRESSOUT_F13_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F13_G);
inv_8850: a_SADDRESSOUT_F13_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8851: a_EQ859 <=  n_10105  XOR n_10115;
or3_8852: n_10105 <=  n_10106  OR n_10109  OR n_10112;
and2_8853: n_10106 <=  n_10107  AND n_10108;
delay_8854: n_10107  <= TRANSPORT a_N1019_aNOT  ;
inv_8855: n_10108  <= TRANSPORT NOT startdma  ;
and2_8856: n_10109 <=  n_10110  AND n_10111;
delay_8857: n_10110  <= TRANSPORT a_LC5_E14  ;
delay_8858: n_10111  <= TRANSPORT startdma  ;
and2_8859: n_10112 <=  n_10113  AND n_10114;
delay_8860: n_10113  <= TRANSPORT a_LC6_E14  ;
delay_8861: n_10114  <= TRANSPORT startdma  ;
and1_8862: n_10115 <=  gnd;
delay_8863: n_10116  <= TRANSPORT clk  ;
filter_8864: FILTER_a8237

    PORT MAP (IN1 => n_10116, Y => a_SADDRESSOUT_F13_G_aCLK);
delay_8865: a_LC7_D6  <= TRANSPORT a_EQ407  ;
xor2_8866: a_EQ407 <=  n_10120  XOR n_10127;
or2_8867: n_10120 <=  n_10121  OR n_10124;
and2_8868: n_10121 <=  n_10122  AND n_10123;
inv_8869: n_10122  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_8870: n_10123  <= TRANSPORT a_SCH0ADDRREG_F15_G  ;
and2_8871: n_10124 <=  n_10125  AND n_10126;
inv_8872: n_10125  <= TRANSPORT NOT a_N2376  ;
delay_8873: n_10126  <= TRANSPORT a_SCH2ADDRREG_F15_G  ;
and1_8874: n_10127 <=  gnd;
delay_8875: a_N1298_aNOT  <= TRANSPORT a_EQ411  ;
xor2_8876: a_EQ411 <=  n_10130  XOR n_10137;
or2_8877: n_10130 <=  n_10131  OR n_10134;
and2_8878: n_10131 <=  n_10132  AND n_10133;
delay_8879: n_10132  <= TRANSPORT a_N2557  ;
delay_8880: n_10133  <= TRANSPORT a_N2555  ;
and2_8881: n_10134 <=  n_10135  AND n_10136;
inv_8882: n_10135  <= TRANSPORT NOT a_N2557  ;
delay_8883: n_10136  <= TRANSPORT a_SADDRESSOUT_F15_G  ;
and1_8884: n_10137 <=  gnd;
delay_8885: a_N1292  <= TRANSPORT a_EQ406  ;
xor2_8886: a_EQ406 <=  n_10140  XOR n_10147;
or2_8887: n_10140 <=  n_10141  OR n_10144;
and2_8888: n_10141 <=  n_10142  AND n_10143;
delay_8889: n_10142  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_8890: n_10143  <= TRANSPORT a_SCH1ADDRREG_F15_G  ;
and2_8891: n_10144 <=  n_10145  AND n_10146;
inv_8892: n_10145  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_8893: n_10146  <= TRANSPORT a_SCH0ADDRREG_F15_G  ;
and1_8894: n_10147 <=  gnd;
delay_8895: a_N1291  <= TRANSPORT a_EQ405  ;
xor2_8896: a_EQ405 <=  n_10150  XOR n_10159;
or3_8897: n_10150 <=  n_10151  OR n_10153  OR n_10156;
and1_8898: n_10151 <=  n_10152;
delay_8899: n_10152  <= TRANSPORT startdma  ;
and2_8900: n_10153 <=  n_10154  AND n_10155;
inv_8901: n_10154  <= TRANSPORT NOT a_N2531  ;
delay_8902: n_10155  <= TRANSPORT a_N1298_aNOT  ;
and2_8903: n_10156 <=  n_10157  AND n_10158;
delay_8904: n_10157  <= TRANSPORT a_N2531  ;
delay_8905: n_10158  <= TRANSPORT a_N1292  ;
and1_8906: n_10159 <=  gnd;
delay_8907: a_LC1_D14  <= TRANSPORT a_EQ408  ;
xor2_8908: a_EQ408 <=  n_10162  XOR n_10169;
or2_8909: n_10162 <=  n_10163  OR n_10166;
and2_8910: n_10163 <=  n_10164  AND n_10165;
inv_8911: n_10164  <= TRANSPORT NOT a_N2377  ;
delay_8912: n_10165  <= TRANSPORT a_SCH3ADDRREG_F15_G  ;
and2_8913: n_10166 <=  n_10167  AND n_10168;
inv_8914: n_10167  <= TRANSPORT NOT a_N88_aNOT  ;
delay_8915: n_10168  <= TRANSPORT a_SCH1ADDRREG_F15_G  ;
and1_8916: n_10169 <=  gnd;
dff_8917: DFF_a8237

    PORT MAP ( D => a_EQ861, CLK => a_SADDRESSOUT_F15_G_aCLK, CLRN => a_SADDRESSOUT_F15_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F15_G);
inv_8918: a_SADDRESSOUT_F15_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8919: a_EQ861 <=  n_10176  XOR n_10186;
or3_8920: n_10176 <=  n_10177  OR n_10180  OR n_10183;
and2_8921: n_10177 <=  n_10178  AND n_10179;
delay_8922: n_10178  <= TRANSPORT a_LC7_D6  ;
delay_8923: n_10179  <= TRANSPORT a_N1291  ;
and2_8924: n_10180 <=  n_10181  AND n_10182;
delay_8925: n_10181  <= TRANSPORT a_N1291  ;
inv_8926: n_10182  <= TRANSPORT NOT startdma  ;
and2_8927: n_10183 <=  n_10184  AND n_10185;
delay_8928: n_10184  <= TRANSPORT a_N1291  ;
delay_8929: n_10185  <= TRANSPORT a_LC1_D14  ;
and1_8930: n_10186 <=  gnd;
delay_8931: n_10187  <= TRANSPORT clk  ;
filter_8932: FILTER_a8237

    PORT MAP (IN1 => n_10187, Y => a_SADDRESSOUT_F15_G_aCLK);
delay_8933: a_SHRQ  <= TRANSPORT a_EQ1132  ;
xor2_8934: a_EQ1132 <=  n_10190  XOR n_10197;
or2_8935: n_10190 <=  n_10191  OR n_10194;
and2_8936: n_10191 <=  n_10192  AND n_10193;
delay_8937: n_10192  <= TRANSPORT a_N2563_aNOT  ;
delay_8938: n_10193  <= TRANSPORT a_N823  ;
and2_8939: n_10194 <=  n_10195  AND n_10196;
delay_8940: n_10195  <= TRANSPORT a_N2563_aNOT  ;
delay_8941: n_10196  <= TRANSPORT a_N1566  ;
and1_8942: n_10197 <=  gnd;
dff_8943: DFF_a8237

    PORT MAP ( D => a_EQ310, CLK => a_N825_aCLK, CLRN => a_N825_aCLRN, PRN => vcc,
          Q => a_N825);
inv_8944: a_N825_aCLRN  <= TRANSPORT NOT reset  ;
xor2_8945: a_EQ310 <=  n_10205  XOR n_10212;
or2_8946: n_10205 <=  n_10206  OR n_10209;
and2_8947: n_10206 <=  n_10207  AND n_10208;
delay_8948: n_10207  <= TRANSPORT a_SHRQ  ;
delay_8949: n_10208  <= TRANSPORT a_N825  ;
and2_8950: n_10209 <=  n_10210  AND n_10211;
delay_8951: n_10210  <= TRANSPORT a_SHRQ  ;
inv_8952: n_10211  <= TRANSPORT NOT neopin  ;
and1_8953: n_10212 <=  gnd;
delay_8954: n_10213  <= TRANSPORT clk  ;
filter_8955: FILTER_a8237

    PORT MAP (IN1 => n_10213, Y => a_N825_aCLK);
delay_8956: a_LC6_E3  <= TRANSPORT a_EQ233  ;
xor2_8957: a_EQ233 <=  n_10217  XOR n_10228;
or3_8958: n_10217 <=  n_10218  OR n_10221  OR n_10224;
and2_8959: n_10218 <=  n_10219  AND n_10220;
inv_8960: n_10219  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
delay_8961: n_10220  <= TRANSPORT a_N3543  ;
and2_8962: n_10221 <=  n_10222  AND n_10223;
inv_8963: n_10222  <= TRANSPORT NOT a_N2557  ;
delay_8964: n_10223  <= TRANSPORT a_N3543  ;
and3_8965: n_10224 <=  n_10225  AND n_10226  AND n_10227;
delay_8966: n_10225  <= TRANSPORT a_N2557  ;
delay_8967: n_10226  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_8968: n_10227  <= TRANSPORT NOT a_N3543  ;
and1_8969: n_10228 <=  gnd;
delay_8970: a_LC4_E3  <= TRANSPORT a_EQ232  ;
xor2_8971: a_EQ232 <=  n_10231  XOR n_10238;
or2_8972: n_10231 <=  n_10232  OR n_10235;
and2_8973: n_10232 <=  n_10233  AND n_10234;
delay_8974: n_10233  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_8975: n_10234  <= TRANSPORT a_SH1WRDCNTREG_F13_G  ;
and2_8976: n_10235 <=  n_10236  AND n_10237;
inv_8977: n_10236  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_8978: n_10237  <= TRANSPORT a_SH0WRDCNTREG_F13_G  ;
and1_8979: n_10238 <=  gnd;
delay_8980: a_N340_aNOT  <= TRANSPORT a_EQ234  ;
xor2_8981: a_EQ234 <=  n_10241  XOR n_10248;
or2_8982: n_10241 <=  n_10242  OR n_10245;
and2_8983: n_10242 <=  n_10243  AND n_10244;
inv_8984: n_10243  <= TRANSPORT NOT a_N2531  ;
delay_8985: n_10244  <= TRANSPORT a_LC6_E3  ;
and2_8986: n_10245 <=  n_10246  AND n_10247;
delay_8987: n_10246  <= TRANSPORT a_N2531  ;
delay_8988: n_10247  <= TRANSPORT a_LC4_E3  ;
and1_8989: n_10248 <=  gnd;
delay_8990: a_LC3_E3  <= TRANSPORT a_EQ231  ;
xor2_8991: a_EQ231 <=  n_10251  XOR n_10258;
or2_8992: n_10251 <=  n_10252  OR n_10255;
and2_8993: n_10252 <=  n_10253  AND n_10254;
inv_8994: n_10253  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_8995: n_10254  <= TRANSPORT a_SH0WRDCNTREG_F13_G  ;
and2_8996: n_10255 <=  n_10256  AND n_10257;
inv_8997: n_10256  <= TRANSPORT NOT a_N2376  ;
delay_8998: n_10257  <= TRANSPORT a_SH2WRDCNTREG_F13_G  ;
and1_8999: n_10258 <=  gnd;
delay_9000: a_LC2_E3  <= TRANSPORT a_EQ230  ;
xor2_9001: a_EQ230 <=  n_10261  XOR n_10268;
or2_9002: n_10261 <=  n_10262  OR n_10265;
and2_9003: n_10262 <=  n_10263  AND n_10264;
inv_9004: n_10263  <= TRANSPORT NOT a_N2377  ;
delay_9005: n_10264  <= TRANSPORT a_SH3WRDCNTREG_F13_G  ;
and2_9006: n_10265 <=  n_10266  AND n_10267;
inv_9007: n_10266  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9008: n_10267  <= TRANSPORT a_SH1WRDCNTREG_F13_G  ;
and1_9009: n_10268 <=  gnd;
dff_9010: DFF_a8237

    PORT MAP ( D => a_EQ839, CLK => a_N3543_aCLK, CLRN => a_N3543_aCLRN, PRN => vcc,
          Q => a_N3543);
inv_9011: a_N3543_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9012: a_EQ839 <=  n_10275  XOR n_10285;
or3_9013: n_10275 <=  n_10276  OR n_10279  OR n_10282;
and2_9014: n_10276 <=  n_10277  AND n_10278;
delay_9015: n_10277  <= TRANSPORT a_N340_aNOT  ;
inv_9016: n_10278  <= TRANSPORT NOT startdma  ;
and2_9017: n_10279 <=  n_10280  AND n_10281;
delay_9018: n_10280  <= TRANSPORT a_LC3_E3  ;
delay_9019: n_10281  <= TRANSPORT startdma  ;
and2_9020: n_10282 <=  n_10283  AND n_10284;
delay_9021: n_10283  <= TRANSPORT a_LC2_E3  ;
delay_9022: n_10284  <= TRANSPORT startdma  ;
and1_9023: n_10285 <=  gnd;
delay_9024: n_10286  <= TRANSPORT clk  ;
filter_9025: FILTER_a8237

    PORT MAP (IN1 => n_10286, Y => a_N3543_aCLK);
delay_9026: a_N866_aNOT  <= TRANSPORT a_EQ317  ;
xor2_9027: a_EQ317 <=  n_10290  XOR n_10305;
or4_9028: n_10290 <=  n_10291  OR n_10294  OR n_10297  OR n_10300;
and2_9029: n_10291 <=  n_10292  AND n_10293;
inv_9030: n_10292  <= TRANSPORT NOT a_LC1_A20_aNOT  ;
delay_9031: n_10293  <= TRANSPORT a_N3542  ;
and2_9032: n_10294 <=  n_10295  AND n_10296;
inv_9033: n_10295  <= TRANSPORT NOT a_N2557  ;
delay_9034: n_10296  <= TRANSPORT a_N3542  ;
and2_9035: n_10297 <=  n_10298  AND n_10299;
delay_9036: n_10298  <= TRANSPORT a_N3543  ;
delay_9037: n_10299  <= TRANSPORT a_N3542  ;
and4_9038: n_10300 <=  n_10301  AND n_10302  AND n_10303  AND n_10304;
delay_9039: n_10301  <= TRANSPORT a_N2557  ;
delay_9040: n_10302  <= TRANSPORT a_LC1_A20_aNOT  ;
inv_9041: n_10303  <= TRANSPORT NOT a_N3543  ;
inv_9042: n_10304  <= TRANSPORT NOT a_N3542  ;
and1_9043: n_10305 <=  gnd;
delay_9044: a_N874  <= TRANSPORT a_EQ321  ;
xor2_9045: a_EQ321 <=  n_10308  XOR n_10315;
or2_9046: n_10308 <=  n_10309  OR n_10312;
and2_9047: n_10309 <=  n_10310  AND n_10311;
inv_9048: n_10310  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9049: n_10311  <= TRANSPORT a_SH0WRDCNTREG_F14_G  ;
and2_9050: n_10312 <=  n_10313  AND n_10314;
delay_9051: n_10313  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9052: n_10314  <= TRANSPORT a_SH1WRDCNTREG_F14_G  ;
and1_9053: n_10315 <=  gnd;
delay_9054: a_LC8_E16  <= TRANSPORT a_EQ322  ;
xor2_9055: a_EQ322 <=  n_10318  XOR n_10325;
or2_9056: n_10318 <=  n_10319  OR n_10322;
and2_9057: n_10319 <=  n_10320  AND n_10321;
inv_9058: n_10320  <= TRANSPORT NOT a_N2531  ;
delay_9059: n_10321  <= TRANSPORT a_N866_aNOT  ;
and2_9060: n_10322 <=  n_10323  AND n_10324;
delay_9061: n_10323  <= TRANSPORT a_N2531  ;
delay_9062: n_10324  <= TRANSPORT a_N874  ;
and1_9063: n_10325 <=  gnd;
delay_9064: a_LC2_E16  <= TRANSPORT a_EQ320  ;
xor2_9065: a_EQ320 <=  n_10328  XOR n_10335;
or2_9066: n_10328 <=  n_10329  OR n_10332;
and2_9067: n_10329 <=  n_10330  AND n_10331;
inv_9068: n_10330  <= TRANSPORT NOT a_N2377  ;
delay_9069: n_10331  <= TRANSPORT a_SH3WRDCNTREG_F14_G  ;
and2_9070: n_10332 <=  n_10333  AND n_10334;
inv_9071: n_10333  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9072: n_10334  <= TRANSPORT a_SH1WRDCNTREG_F14_G  ;
and1_9073: n_10335 <=  gnd;
delay_9074: a_LC1_E16  <= TRANSPORT a_EQ319  ;
xor2_9075: a_EQ319 <=  n_10338  XOR n_10345;
or2_9076: n_10338 <=  n_10339  OR n_10342;
and2_9077: n_10339 <=  n_10340  AND n_10341;
inv_9078: n_10340  <= TRANSPORT NOT a_N2376  ;
delay_9079: n_10341  <= TRANSPORT a_SH2WRDCNTREG_F14_G  ;
and2_9080: n_10342 <=  n_10343  AND n_10344;
inv_9081: n_10343  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9082: n_10344  <= TRANSPORT a_SH0WRDCNTREG_F14_G  ;
and1_9083: n_10345 <=  gnd;
dff_9084: DFF_a8237

    PORT MAP ( D => a_EQ838, CLK => a_N3542_aCLK, CLRN => a_N3542_aCLRN, PRN => vcc,
          Q => a_N3542);
inv_9085: a_N3542_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9086: a_EQ838 <=  n_10352  XOR n_10362;
or3_9087: n_10352 <=  n_10353  OR n_10356  OR n_10359;
and2_9088: n_10353 <=  n_10354  AND n_10355;
delay_9089: n_10354  <= TRANSPORT a_LC8_E16  ;
inv_9090: n_10355  <= TRANSPORT NOT startdma  ;
and2_9091: n_10356 <=  n_10357  AND n_10358;
delay_9092: n_10357  <= TRANSPORT a_LC2_E16  ;
delay_9093: n_10358  <= TRANSPORT startdma  ;
and2_9094: n_10359 <=  n_10360  AND n_10361;
delay_9095: n_10360  <= TRANSPORT a_LC1_E16  ;
delay_9096: n_10361  <= TRANSPORT startdma  ;
and1_9097: n_10362 <=  gnd;
delay_9098: n_10363  <= TRANSPORT clk  ;
filter_9099: FILTER_a8237

    PORT MAP (IN1 => n_10363, Y => a_N3542_aCLK);
delay_9100: a_N2372_aNOT  <= TRANSPORT a_N2372_aNOT_aIN  ;
xor2_9101: a_N2372_aNOT_aIN <=  n_10367  XOR n_10373;
or1_9102: n_10367 <=  n_10368;
and4_9103: n_10368 <=  n_10369  AND n_10370  AND n_10371  AND n_10372;
delay_9104: n_10369  <= TRANSPORT a_N820  ;
inv_9105: n_10370  <= TRANSPORT NOT a_N822  ;
inv_9106: n_10371  <= TRANSPORT NOT a_N821  ;
delay_9107: n_10372  <= TRANSPORT a_N823  ;
and1_9108: n_10373 <=  gnd;
dff_9109: DFF_a8237

    PORT MAP ( D => a_EQ1181, CLK => a_STEMPORARYREG_F0_G_aCLK, CLRN => a_STEMPORARYREG_F0_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F0_G);
inv_9110: a_STEMPORARYREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9111: a_EQ1181 <=  n_10381  XOR n_10390;
or2_9112: n_10381 <=  n_10382  OR n_10386;
and3_9113: n_10382 <=  n_10383  AND n_10384  AND n_10385;
delay_9114: n_10383  <= TRANSPORT a_N2563_aNOT  ;
inv_9115: n_10384  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9116: n_10385  <= TRANSPORT a_STEMPORARYREG_F0_G  ;
and3_9117: n_10386 <=  n_10387  AND n_10388  AND n_10389;
delay_9118: n_10387  <= TRANSPORT a_N2563_aNOT  ;
delay_9119: n_10388  <= TRANSPORT dbin(0)  ;
delay_9120: n_10389  <= TRANSPORT a_N2372_aNOT  ;
and1_9121: n_10390 <=  gnd;
delay_9122: n_10391  <= TRANSPORT clk  ;
filter_9123: FILTER_a8237

    PORT MAP (IN1 => n_10391, Y => a_STEMPORARYREG_F0_G_aCLK);
delay_9124: a_N1338_aNOT  <= TRANSPORT a_EQ425  ;
xor2_9125: a_EQ425 <=  n_10395  XOR n_10402;
or2_9126: n_10395 <=  n_10396  OR n_10399;
and2_9127: n_10396 <=  n_10397  AND n_10398;
delay_9128: n_10397  <= TRANSPORT a_N2557  ;
delay_9129: n_10398  <= TRANSPORT a_N2548  ;
and2_9130: n_10399 <=  n_10400  AND n_10401;
inv_9131: n_10400  <= TRANSPORT NOT a_N2557  ;
delay_9132: n_10401  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and1_9133: n_10402 <=  gnd;
delay_9134: a_N1327  <= TRANSPORT a_EQ417  ;
xor2_9135: a_EQ417 <=  n_10405  XOR n_10412;
or2_9136: n_10405 <=  n_10406  OR n_10409;
and2_9137: n_10406 <=  n_10407  AND n_10408;
inv_9138: n_10407  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9139: n_10408  <= TRANSPORT a_SCH0ADDRREG_F8_G  ;
and2_9140: n_10409 <=  n_10410  AND n_10411;
delay_9141: n_10410  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9142: n_10411  <= TRANSPORT a_SCH1ADDRREG_F8_G  ;
and1_9143: n_10412 <=  gnd;
delay_9144: a_LC6_F5  <= TRANSPORT a_EQ416  ;
xor2_9145: a_EQ416 <=  n_10415  XOR n_10422;
or2_9146: n_10415 <=  n_10416  OR n_10419;
and2_9147: n_10416 <=  n_10417  AND n_10418;
inv_9148: n_10417  <= TRANSPORT NOT a_N2531  ;
delay_9149: n_10418  <= TRANSPORT a_N1338_aNOT  ;
and2_9150: n_10419 <=  n_10420  AND n_10421;
delay_9151: n_10420  <= TRANSPORT a_N2531  ;
delay_9152: n_10421  <= TRANSPORT a_N1327  ;
and1_9153: n_10422 <=  gnd;
delay_9154: a_LC1_F5  <= TRANSPORT a_EQ419  ;
xor2_9155: a_EQ419 <=  n_10425  XOR n_10432;
or2_9156: n_10425 <=  n_10426  OR n_10429;
and2_9157: n_10426 <=  n_10427  AND n_10428;
inv_9158: n_10427  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9159: n_10428  <= TRANSPORT a_SCH1ADDRREG_F8_G  ;
and2_9160: n_10429 <=  n_10430  AND n_10431;
inv_9161: n_10430  <= TRANSPORT NOT a_N2377  ;
delay_9162: n_10431  <= TRANSPORT a_SCH3ADDRREG_F8_G  ;
and1_9163: n_10432 <=  gnd;
delay_9164: a_LC2_F5  <= TRANSPORT a_EQ418  ;
xor2_9165: a_EQ418 <=  n_10435  XOR n_10442;
or2_9166: n_10435 <=  n_10436  OR n_10439;
and2_9167: n_10436 <=  n_10437  AND n_10438;
inv_9168: n_10437  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9169: n_10438  <= TRANSPORT a_SCH0ADDRREG_F8_G  ;
and2_9170: n_10439 <=  n_10440  AND n_10441;
inv_9171: n_10440  <= TRANSPORT NOT a_N2376  ;
delay_9172: n_10441  <= TRANSPORT a_SCH2ADDRREG_F8_G  ;
and1_9173: n_10442 <=  gnd;
dff_9174: DFF_a8237

    PORT MAP ( D => a_EQ854, CLK => a_SADDRESSOUT_F8_G_aCLK, CLRN => a_SADDRESSOUT_F8_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F8_G);
inv_9175: a_SADDRESSOUT_F8_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9176: a_EQ854 <=  n_10449  XOR n_10459;
or3_9177: n_10449 <=  n_10450  OR n_10453  OR n_10456;
and2_9178: n_10450 <=  n_10451  AND n_10452;
delay_9179: n_10451  <= TRANSPORT a_LC6_F5  ;
inv_9180: n_10452  <= TRANSPORT NOT startdma  ;
and2_9181: n_10453 <=  n_10454  AND n_10455;
delay_9182: n_10454  <= TRANSPORT a_LC1_F5  ;
delay_9183: n_10455  <= TRANSPORT startdma  ;
and2_9184: n_10456 <=  n_10457  AND n_10458;
delay_9185: n_10457  <= TRANSPORT a_LC2_F5  ;
delay_9186: n_10458  <= TRANSPORT startdma  ;
and1_9187: n_10459 <=  gnd;
delay_9188: n_10460  <= TRANSPORT clk  ;
filter_9189: FILTER_a8237

    PORT MAP (IN1 => n_10460, Y => a_SADDRESSOUT_F8_G_aCLK);
dff_9190: DFF_a8237

    PORT MAP ( D => a_EQ1123, CLK => a_SCOMMANDREG_F0_G_aCLK, CLRN => a_SCOMMANDREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F0_G);
inv_9191: a_SCOMMANDREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9192: a_EQ1123 <=  n_10468  XOR n_10477;
or2_9193: n_10468 <=  n_10469  OR n_10473;
and3_9194: n_10469 <=  n_10470  AND n_10471  AND n_10472;
delay_9195: n_10470  <= TRANSPORT a_N2563_aNOT  ;
delay_9196: n_10471  <= TRANSPORT a_N2571_aNOT  ;
delay_9197: n_10472  <= TRANSPORT a_SCOMMANDREG_F0_G  ;
and3_9198: n_10473 <=  n_10474  AND n_10475  AND n_10476;
delay_9199: n_10474  <= TRANSPORT a_N2563_aNOT  ;
delay_9200: n_10475  <= TRANSPORT dbin(0)  ;
inv_9201: n_10476  <= TRANSPORT NOT a_N2571_aNOT  ;
and1_9202: n_10477 <=  gnd;
delay_9203: n_10478  <= TRANSPORT clk  ;
filter_9204: FILTER_a8237

    PORT MAP (IN1 => n_10478, Y => a_SCOMMANDREG_F0_G_aCLK);
dff_9205: DFF_a8237

    PORT MAP ( D => a_EQ1182, CLK => a_STEMPORARYREG_F1_G_aCLK, CLRN => a_STEMPORARYREG_F1_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F1_G);
inv_9206: a_STEMPORARYREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9207: a_EQ1182 <=  n_10487  XOR n_10496;
or2_9208: n_10487 <=  n_10488  OR n_10492;
and3_9209: n_10488 <=  n_10489  AND n_10490  AND n_10491;
delay_9210: n_10489  <= TRANSPORT a_N2563_aNOT  ;
inv_9211: n_10490  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9212: n_10491  <= TRANSPORT a_STEMPORARYREG_F1_G  ;
and3_9213: n_10492 <=  n_10493  AND n_10494  AND n_10495;
delay_9214: n_10493  <= TRANSPORT a_N2563_aNOT  ;
delay_9215: n_10494  <= TRANSPORT dbin(1)  ;
delay_9216: n_10495  <= TRANSPORT a_N2372_aNOT  ;
and1_9217: n_10496 <=  gnd;
delay_9218: n_10497  <= TRANSPORT clk  ;
filter_9219: FILTER_a8237

    PORT MAP (IN1 => n_10497, Y => a_STEMPORARYREG_F1_G_aCLK);
delay_9220: a_LC2_A18  <= TRANSPORT a_EQ279  ;
xor2_9221: a_EQ279 <=  n_10501  XOR n_10508;
or2_9222: n_10501 <=  n_10502  OR n_10505;
and2_9223: n_10502 <=  n_10503  AND n_10504;
delay_9224: n_10503  <= TRANSPORT a_N2557  ;
delay_9225: n_10504  <= TRANSPORT a_N2549  ;
and2_9226: n_10505 <=  n_10506  AND n_10507;
inv_9227: n_10506  <= TRANSPORT NOT a_N2557  ;
delay_9228: n_10507  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
and1_9229: n_10508 <=  gnd;
delay_9230: a_LC1_A18  <= TRANSPORT a_EQ280  ;
xor2_9231: a_EQ280 <=  n_10511  XOR n_10518;
or2_9232: n_10511 <=  n_10512  OR n_10515;
and2_9233: n_10512 <=  n_10513  AND n_10514;
delay_9234: n_10513  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9235: n_10514  <= TRANSPORT a_SCH1ADDRREG_F9_G  ;
and2_9236: n_10515 <=  n_10516  AND n_10517;
inv_9237: n_10516  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9238: n_10517  <= TRANSPORT a_SCH0ADDRREG_F9_G  ;
and1_9239: n_10518 <=  gnd;
delay_9240: a_N672_aNOT  <= TRANSPORT a_EQ283  ;
xor2_9241: a_EQ283 <=  n_10521  XOR n_10528;
or2_9242: n_10521 <=  n_10522  OR n_10525;
and2_9243: n_10522 <=  n_10523  AND n_10524;
inv_9244: n_10523  <= TRANSPORT NOT a_N2531  ;
delay_9245: n_10524  <= TRANSPORT a_LC2_A18  ;
and2_9246: n_10525 <=  n_10526  AND n_10527;
delay_9247: n_10526  <= TRANSPORT a_N2531  ;
delay_9248: n_10527  <= TRANSPORT a_LC1_A18  ;
and1_9249: n_10528 <=  gnd;
delay_9250: a_LC4_A18  <= TRANSPORT a_EQ282  ;
xor2_9251: a_EQ282 <=  n_10531  XOR n_10538;
or2_9252: n_10531 <=  n_10532  OR n_10535;
and2_9253: n_10532 <=  n_10533  AND n_10534;
inv_9254: n_10533  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9255: n_10534  <= TRANSPORT a_SCH1ADDRREG_F9_G  ;
and2_9256: n_10535 <=  n_10536  AND n_10537;
inv_9257: n_10536  <= TRANSPORT NOT a_N2377  ;
delay_9258: n_10537  <= TRANSPORT a_SCH3ADDRREG_F9_G  ;
and1_9259: n_10538 <=  gnd;
delay_9260: a_LC5_A18  <= TRANSPORT a_EQ281  ;
xor2_9261: a_EQ281 <=  n_10541  XOR n_10548;
or2_9262: n_10541 <=  n_10542  OR n_10545;
and2_9263: n_10542 <=  n_10543  AND n_10544;
inv_9264: n_10543  <= TRANSPORT NOT a_N2376  ;
delay_9265: n_10544  <= TRANSPORT a_SCH2ADDRREG_F9_G  ;
and2_9266: n_10545 <=  n_10546  AND n_10547;
inv_9267: n_10546  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9268: n_10547  <= TRANSPORT a_SCH0ADDRREG_F9_G  ;
and1_9269: n_10548 <=  gnd;
dff_9270: DFF_a8237

    PORT MAP ( D => a_EQ855, CLK => a_SADDRESSOUT_F9_G_aCLK, CLRN => a_SADDRESSOUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F9_G);
inv_9271: a_SADDRESSOUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9272: a_EQ855 <=  n_10555  XOR n_10565;
or3_9273: n_10555 <=  n_10556  OR n_10559  OR n_10562;
and2_9274: n_10556 <=  n_10557  AND n_10558;
delay_9275: n_10557  <= TRANSPORT a_N672_aNOT  ;
inv_9276: n_10558  <= TRANSPORT NOT startdma  ;
and2_9277: n_10559 <=  n_10560  AND n_10561;
delay_9278: n_10560  <= TRANSPORT a_LC4_A18  ;
delay_9279: n_10561  <= TRANSPORT startdma  ;
and2_9280: n_10562 <=  n_10563  AND n_10564;
delay_9281: n_10563  <= TRANSPORT a_LC5_A18  ;
delay_9282: n_10564  <= TRANSPORT startdma  ;
and1_9283: n_10565 <=  gnd;
delay_9284: n_10566  <= TRANSPORT clk  ;
filter_9285: FILTER_a8237

    PORT MAP (IN1 => n_10566, Y => a_SADDRESSOUT_F9_G_aCLK);
delay_9286: a_LC3_E15  <= TRANSPORT a_EQ333  ;
xor2_9287: a_EQ333 <=  n_10570  XOR n_10577;
or2_9288: n_10570 <=  n_10571  OR n_10574;
and2_9289: n_10571 <=  n_10572  AND n_10573;
delay_9290: n_10572  <= TRANSPORT a_N2557  ;
delay_9291: n_10573  <= TRANSPORT a_N2550  ;
and2_9292: n_10574 <=  n_10575  AND n_10576;
inv_9293: n_10575  <= TRANSPORT NOT a_N2557  ;
delay_9294: n_10576  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and1_9295: n_10577 <=  gnd;
delay_9296: a_LC1_E18  <= TRANSPORT a_EQ332  ;
xor2_9297: a_EQ332 <=  n_10580  XOR n_10587;
or2_9298: n_10580 <=  n_10581  OR n_10584;
and2_9299: n_10581 <=  n_10582  AND n_10583;
delay_9300: n_10582  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9301: n_10583  <= TRANSPORT a_SCH1ADDRREG_F10_G  ;
and2_9302: n_10584 <=  n_10585  AND n_10586;
inv_9303: n_10585  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9304: n_10586  <= TRANSPORT a_SCH0ADDRREG_F10_G  ;
and1_9305: n_10587 <=  gnd;
delay_9306: a_N1000_aNOT  <= TRANSPORT a_EQ336  ;
xor2_9307: a_EQ336 <=  n_10590  XOR n_10597;
or2_9308: n_10590 <=  n_10591  OR n_10594;
and2_9309: n_10591 <=  n_10592  AND n_10593;
inv_9310: n_10592  <= TRANSPORT NOT a_N2531  ;
delay_9311: n_10593  <= TRANSPORT a_LC3_E15  ;
and2_9312: n_10594 <=  n_10595  AND n_10596;
delay_9313: n_10595  <= TRANSPORT a_N2531  ;
delay_9314: n_10596  <= TRANSPORT a_LC1_E18  ;
and1_9315: n_10597 <=  gnd;
delay_9316: a_LC1_E21  <= TRANSPORT a_EQ335  ;
xor2_9317: a_EQ335 <=  n_10600  XOR n_10607;
or2_9318: n_10600 <=  n_10601  OR n_10604;
and2_9319: n_10601 <=  n_10602  AND n_10603;
inv_9320: n_10602  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9321: n_10603  <= TRANSPORT a_SCH0ADDRREG_F10_G  ;
and2_9322: n_10604 <=  n_10605  AND n_10606;
inv_9323: n_10605  <= TRANSPORT NOT a_N2376  ;
delay_9324: n_10606  <= TRANSPORT a_SCH2ADDRREG_F10_G  ;
and1_9325: n_10607 <=  gnd;
delay_9326: a_LC8_E15  <= TRANSPORT a_EQ334  ;
xor2_9327: a_EQ334 <=  n_10610  XOR n_10617;
or2_9328: n_10610 <=  n_10611  OR n_10614;
and2_9329: n_10611 <=  n_10612  AND n_10613;
inv_9330: n_10612  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9331: n_10613  <= TRANSPORT a_SCH1ADDRREG_F10_G  ;
and2_9332: n_10614 <=  n_10615  AND n_10616;
inv_9333: n_10615  <= TRANSPORT NOT a_N2377  ;
delay_9334: n_10616  <= TRANSPORT a_SCH3ADDRREG_F10_G  ;
and1_9335: n_10617 <=  gnd;
dff_9336: DFF_a8237

    PORT MAP ( D => a_EQ856, CLK => a_SADDRESSOUT_F10_G_aCLK, CLRN => a_SADDRESSOUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F10_G);
inv_9337: a_SADDRESSOUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9338: a_EQ856 <=  n_10624  XOR n_10634;
or3_9339: n_10624 <=  n_10625  OR n_10628  OR n_10631;
and2_9340: n_10625 <=  n_10626  AND n_10627;
delay_9341: n_10626  <= TRANSPORT a_N1000_aNOT  ;
inv_9342: n_10627  <= TRANSPORT NOT startdma  ;
and2_9343: n_10628 <=  n_10629  AND n_10630;
delay_9344: n_10629  <= TRANSPORT a_LC1_E21  ;
delay_9345: n_10630  <= TRANSPORT startdma  ;
and2_9346: n_10631 <=  n_10632  AND n_10633;
delay_9347: n_10632  <= TRANSPORT a_LC8_E15  ;
delay_9348: n_10633  <= TRANSPORT startdma  ;
and1_9349: n_10634 <=  gnd;
delay_9350: n_10635  <= TRANSPORT clk  ;
filter_9351: FILTER_a8237

    PORT MAP (IN1 => n_10635, Y => a_SADDRESSOUT_F10_G_aCLK);
dff_9352: DFF_a8237

    PORT MAP ( D => a_EQ1183, CLK => a_STEMPORARYREG_F2_G_aCLK, CLRN => a_STEMPORARYREG_F2_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F2_G);
inv_9353: a_STEMPORARYREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9354: a_EQ1183 <=  n_10644  XOR n_10653;
or2_9355: n_10644 <=  n_10645  OR n_10649;
and3_9356: n_10645 <=  n_10646  AND n_10647  AND n_10648;
delay_9357: n_10646  <= TRANSPORT a_N2563_aNOT  ;
inv_9358: n_10647  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9359: n_10648  <= TRANSPORT a_STEMPORARYREG_F2_G  ;
and3_9360: n_10649 <=  n_10650  AND n_10651  AND n_10652;
delay_9361: n_10650  <= TRANSPORT a_N2563_aNOT  ;
delay_9362: n_10651  <= TRANSPORT dbin(2)  ;
delay_9363: n_10652  <= TRANSPORT a_N2372_aNOT  ;
and1_9364: n_10653 <=  gnd;
delay_9365: n_10654  <= TRANSPORT clk  ;
filter_9366: FILTER_a8237

    PORT MAP (IN1 => n_10654, Y => a_STEMPORARYREG_F2_G_aCLK);
delay_9367: a_N1339_aNOT  <= TRANSPORT a_EQ426  ;
xor2_9368: a_EQ426 <=  n_10658  XOR n_10665;
or2_9369: n_10658 <=  n_10659  OR n_10662;
and2_9370: n_10659 <=  n_10660  AND n_10661;
delay_9371: n_10660  <= TRANSPORT a_N2557  ;
delay_9372: n_10661  <= TRANSPORT a_N2551  ;
and2_9373: n_10662 <=  n_10663  AND n_10664;
inv_9374: n_10663  <= TRANSPORT NOT a_N2557  ;
delay_9375: n_10664  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and1_9376: n_10665 <=  gnd;
delay_9377: a_N1333  <= TRANSPORT a_EQ421  ;
xor2_9378: a_EQ421 <=  n_10668  XOR n_10675;
or2_9379: n_10668 <=  n_10669  OR n_10672;
and2_9380: n_10669 <=  n_10670  AND n_10671;
delay_9381: n_10670  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9382: n_10671  <= TRANSPORT a_SCH1ADDRREG_F11_G  ;
and2_9383: n_10672 <=  n_10673  AND n_10674;
inv_9384: n_10673  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9385: n_10674  <= TRANSPORT a_SCH0ADDRREG_F11_G  ;
and1_9386: n_10675 <=  gnd;
delay_9387: a_LC3_A19  <= TRANSPORT a_EQ420  ;
xor2_9388: a_EQ420 <=  n_10678  XOR n_10685;
or2_9389: n_10678 <=  n_10679  OR n_10682;
and2_9390: n_10679 <=  n_10680  AND n_10681;
inv_9391: n_10680  <= TRANSPORT NOT a_N2531  ;
delay_9392: n_10681  <= TRANSPORT a_N1339_aNOT  ;
and2_9393: n_10682 <=  n_10683  AND n_10684;
delay_9394: n_10683  <= TRANSPORT a_N2531  ;
delay_9395: n_10684  <= TRANSPORT a_N1333  ;
and1_9396: n_10685 <=  gnd;
delay_9397: a_LC1_A19  <= TRANSPORT a_EQ423  ;
xor2_9398: a_EQ423 <=  n_10688  XOR n_10695;
or2_9399: n_10688 <=  n_10689  OR n_10692;
and2_9400: n_10689 <=  n_10690  AND n_10691;
inv_9401: n_10690  <= TRANSPORT NOT a_N2376  ;
delay_9402: n_10691  <= TRANSPORT a_SCH2ADDRREG_F11_G  ;
and2_9403: n_10692 <=  n_10693  AND n_10694;
inv_9404: n_10693  <= TRANSPORT NOT a_N2377  ;
delay_9405: n_10694  <= TRANSPORT a_SCH3ADDRREG_F11_G  ;
and1_9406: n_10695 <=  gnd;
delay_9407: a_LC2_A19  <= TRANSPORT a_EQ422  ;
xor2_9408: a_EQ422 <=  n_10698  XOR n_10705;
or2_9409: n_10698 <=  n_10699  OR n_10702;
and2_9410: n_10699 <=  n_10700  AND n_10701;
inv_9411: n_10700  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9412: n_10701  <= TRANSPORT a_SCH0ADDRREG_F11_G  ;
and2_9413: n_10702 <=  n_10703  AND n_10704;
inv_9414: n_10703  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9415: n_10704  <= TRANSPORT a_SCH1ADDRREG_F11_G  ;
and1_9416: n_10705 <=  gnd;
dff_9417: DFF_a8237

    PORT MAP ( D => a_EQ857, CLK => a_SADDRESSOUT_F11_G_aCLK, CLRN => a_SADDRESSOUT_F11_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F11_G);
inv_9418: a_SADDRESSOUT_F11_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9419: a_EQ857 <=  n_10712  XOR n_10722;
or3_9420: n_10712 <=  n_10713  OR n_10716  OR n_10719;
and2_9421: n_10713 <=  n_10714  AND n_10715;
delay_9422: n_10714  <= TRANSPORT a_LC3_A19  ;
inv_9423: n_10715  <= TRANSPORT NOT startdma  ;
and2_9424: n_10716 <=  n_10717  AND n_10718;
delay_9425: n_10717  <= TRANSPORT a_LC1_A19  ;
delay_9426: n_10718  <= TRANSPORT startdma  ;
and2_9427: n_10719 <=  n_10720  AND n_10721;
delay_9428: n_10720  <= TRANSPORT a_LC2_A19  ;
delay_9429: n_10721  <= TRANSPORT startdma  ;
and1_9430: n_10722 <=  gnd;
delay_9431: n_10723  <= TRANSPORT clk  ;
filter_9432: FILTER_a8237

    PORT MAP (IN1 => n_10723, Y => a_SADDRESSOUT_F11_G_aCLK);
dff_9433: DFF_a8237

    PORT MAP ( D => a_EQ1184, CLK => a_STEMPORARYREG_F3_G_aCLK, CLRN => a_STEMPORARYREG_F3_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F3_G);
inv_9434: a_STEMPORARYREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9435: a_EQ1184 <=  n_10732  XOR n_10741;
or2_9436: n_10732 <=  n_10733  OR n_10737;
and3_9437: n_10733 <=  n_10734  AND n_10735  AND n_10736;
delay_9438: n_10734  <= TRANSPORT a_N2563_aNOT  ;
inv_9439: n_10735  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9440: n_10736  <= TRANSPORT a_STEMPORARYREG_F3_G  ;
and3_9441: n_10737 <=  n_10738  AND n_10739  AND n_10740;
delay_9442: n_10738  <= TRANSPORT a_N2563_aNOT  ;
delay_9443: n_10739  <= TRANSPORT dbin(3)  ;
delay_9444: n_10740  <= TRANSPORT a_N2372_aNOT  ;
and1_9445: n_10741 <=  gnd;
delay_9446: n_10742  <= TRANSPORT clk  ;
filter_9447: FILTER_a8237

    PORT MAP (IN1 => n_10742, Y => a_STEMPORARYREG_F3_G_aCLK);
delay_9448: a_LC3_A26  <= TRANSPORT a_EQ207  ;
xor2_9449: a_EQ207 <=  n_10746  XOR n_10753;
or2_9450: n_10746 <=  n_10747  OR n_10750;
and2_9451: n_10747 <=  n_10748  AND n_10749;
delay_9452: n_10748  <= TRANSPORT a_N2557  ;
delay_9453: n_10749  <= TRANSPORT a_N2552  ;
and2_9454: n_10750 <=  n_10751  AND n_10752;
inv_9455: n_10751  <= TRANSPORT NOT a_N2557  ;
delay_9456: n_10752  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and1_9457: n_10753 <=  gnd;
delay_9458: a_LC2_A26  <= TRANSPORT a_EQ206  ;
xor2_9459: a_EQ206 <=  n_10756  XOR n_10763;
or2_9460: n_10756 <=  n_10757  OR n_10760;
and2_9461: n_10757 <=  n_10758  AND n_10759;
inv_9462: n_10758  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9463: n_10759  <= TRANSPORT a_SCH0ADDRREG_F12_G  ;
and2_9464: n_10760 <=  n_10761  AND n_10762;
delay_9465: n_10761  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9466: n_10762  <= TRANSPORT a_SCH1ADDRREG_F12_G  ;
and1_9467: n_10763 <=  gnd;
delay_9468: a_LC4_A26  <= TRANSPORT a_EQ210  ;
xor2_9469: a_EQ210 <=  n_10766  XOR n_10773;
or2_9470: n_10766 <=  n_10767  OR n_10770;
and2_9471: n_10767 <=  n_10768  AND n_10769;
inv_9472: n_10768  <= TRANSPORT NOT a_N2531  ;
delay_9473: n_10769  <= TRANSPORT a_LC3_A26  ;
and2_9474: n_10770 <=  n_10771  AND n_10772;
delay_9475: n_10771  <= TRANSPORT a_N2531  ;
delay_9476: n_10772  <= TRANSPORT a_LC2_A26  ;
and1_9477: n_10773 <=  gnd;
delay_9478: a_LC5_A26  <= TRANSPORT a_EQ209  ;
xor2_9479: a_EQ209 <=  n_10776  XOR n_10783;
or2_9480: n_10776 <=  n_10777  OR n_10780;
and2_9481: n_10777 <=  n_10778  AND n_10779;
inv_9482: n_10778  <= TRANSPORT NOT a_N2376  ;
delay_9483: n_10779  <= TRANSPORT a_SCH2ADDRREG_F12_G  ;
and2_9484: n_10780 <=  n_10781  AND n_10782;
inv_9485: n_10781  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9486: n_10782  <= TRANSPORT a_SCH0ADDRREG_F12_G  ;
and1_9487: n_10783 <=  gnd;
delay_9488: a_LC6_A26  <= TRANSPORT a_EQ208  ;
xor2_9489: a_EQ208 <=  n_10786  XOR n_10793;
or2_9490: n_10786 <=  n_10787  OR n_10790;
and2_9491: n_10787 <=  n_10788  AND n_10789;
inv_9492: n_10788  <= TRANSPORT NOT a_N2377  ;
delay_9493: n_10789  <= TRANSPORT a_SCH3ADDRREG_F12_G  ;
and2_9494: n_10790 <=  n_10791  AND n_10792;
inv_9495: n_10791  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9496: n_10792  <= TRANSPORT a_SCH1ADDRREG_F12_G  ;
and1_9497: n_10793 <=  gnd;
dff_9498: DFF_a8237

    PORT MAP ( D => a_EQ858, CLK => a_SADDRESSOUT_F12_G_aCLK, CLRN => a_SADDRESSOUT_F12_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F12_G);
inv_9499: a_SADDRESSOUT_F12_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9500: a_EQ858 <=  n_10800  XOR n_10810;
or3_9501: n_10800 <=  n_10801  OR n_10804  OR n_10807;
and2_9502: n_10801 <=  n_10802  AND n_10803;
delay_9503: n_10802  <= TRANSPORT a_LC4_A26  ;
inv_9504: n_10803  <= TRANSPORT NOT startdma  ;
and2_9505: n_10804 <=  n_10805  AND n_10806;
delay_9506: n_10805  <= TRANSPORT a_LC5_A26  ;
delay_9507: n_10806  <= TRANSPORT startdma  ;
and2_9508: n_10807 <=  n_10808  AND n_10809;
delay_9509: n_10808  <= TRANSPORT a_LC6_A26  ;
delay_9510: n_10809  <= TRANSPORT startdma  ;
and1_9511: n_10810 <=  gnd;
delay_9512: n_10811  <= TRANSPORT clk  ;
filter_9513: FILTER_a8237

    PORT MAP (IN1 => n_10811, Y => a_SADDRESSOUT_F12_G_aCLK);
dff_9514: DFF_a8237

    PORT MAP ( D => a_EQ1129, CLK => a_SCOMMANDREG_F6_G_aCLK, CLRN => a_SCOMMANDREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F6_G);
inv_9515: a_SCOMMANDREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9516: a_EQ1129 <=  n_10820  XOR n_10828;
or2_9517: n_10820 <=  n_10821  OR n_10825;
and3_9518: n_10821 <=  n_10822  AND n_10823  AND n_10824;
delay_9519: n_10822  <= TRANSPORT a_N2563_aNOT  ;
delay_9520: n_10823  <= TRANSPORT a_N2571_aNOT  ;
delay_9521: n_10824  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
and2_9522: n_10825 <=  n_10826  AND n_10827;
inv_9523: n_10826  <= TRANSPORT NOT a_N2571_aNOT  ;
delay_9524: n_10827  <= TRANSPORT dbin(6)  ;
and1_9525: n_10828 <=  gnd;
delay_9526: n_10829  <= TRANSPORT clk  ;
filter_9527: FILTER_a8237

    PORT MAP (IN1 => n_10829, Y => a_SCOMMANDREG_F6_G_aCLK);
dff_9528: DFF_a8237

    PORT MAP ( D => a_EQ1186, CLK => a_STEMPORARYREG_F5_G_aCLK, CLRN => a_STEMPORARYREG_F5_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F5_G);
inv_9529: a_STEMPORARYREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9530: a_EQ1186 <=  n_10838  XOR n_10847;
or2_9531: n_10838 <=  n_10839  OR n_10843;
and3_9532: n_10839 <=  n_10840  AND n_10841  AND n_10842;
delay_9533: n_10840  <= TRANSPORT a_N2563_aNOT  ;
inv_9534: n_10841  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9535: n_10842  <= TRANSPORT a_STEMPORARYREG_F5_G  ;
and3_9536: n_10843 <=  n_10844  AND n_10845  AND n_10846;
delay_9537: n_10844  <= TRANSPORT a_N2563_aNOT  ;
delay_9538: n_10845  <= TRANSPORT a_N2372_aNOT  ;
delay_9539: n_10846  <= TRANSPORT dbin(5)  ;
and1_9540: n_10847 <=  gnd;
delay_9541: n_10848  <= TRANSPORT clk  ;
filter_9542: FILTER_a8237

    PORT MAP (IN1 => n_10848, Y => a_STEMPORARYREG_F5_G_aCLK);
dff_9543: DFF_a8237

    PORT MAP ( D => a_EQ1187, CLK => a_STEMPORARYREG_F6_G_aCLK, CLRN => a_STEMPORARYREG_F6_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F6_G);
inv_9544: a_STEMPORARYREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9545: a_EQ1187 <=  n_10857  XOR n_10866;
or2_9546: n_10857 <=  n_10858  OR n_10862;
and3_9547: n_10858 <=  n_10859  AND n_10860  AND n_10861;
delay_9548: n_10859  <= TRANSPORT a_N2563_aNOT  ;
inv_9549: n_10860  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9550: n_10861  <= TRANSPORT a_STEMPORARYREG_F6_G  ;
and3_9551: n_10862 <=  n_10863  AND n_10864  AND n_10865;
delay_9552: n_10863  <= TRANSPORT a_N2563_aNOT  ;
delay_9553: n_10864  <= TRANSPORT dbin(6)  ;
delay_9554: n_10865  <= TRANSPORT a_N2372_aNOT  ;
and1_9555: n_10866 <=  gnd;
delay_9556: n_10867  <= TRANSPORT clk  ;
filter_9557: FILTER_a8237

    PORT MAP (IN1 => n_10867, Y => a_STEMPORARYREG_F6_G_aCLK);
delay_9558: a_LC4_F9  <= TRANSPORT a_EQ218  ;
xor2_9559: a_EQ218 <=  n_10871  XOR n_10878;
or2_9560: n_10871 <=  n_10872  OR n_10875;
and2_9561: n_10872 <=  n_10873  AND n_10874;
delay_9562: n_10873  <= TRANSPORT a_N2557  ;
delay_9563: n_10874  <= TRANSPORT a_N2554  ;
and2_9564: n_10875 <=  n_10876  AND n_10877;
inv_9565: n_10876  <= TRANSPORT NOT a_N2557  ;
delay_9566: n_10877  <= TRANSPORT a_SADDRESSOUT_F14_G  ;
and1_9567: n_10878 <=  gnd;
delay_9568: a_LC7_F9  <= TRANSPORT a_EQ217  ;
xor2_9569: a_EQ217 <=  n_10881  XOR n_10888;
or2_9570: n_10881 <=  n_10882  OR n_10885;
and2_9571: n_10882 <=  n_10883  AND n_10884;
delay_9572: n_10883  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_9573: n_10884  <= TRANSPORT a_SCH1ADDRREG_F14_G  ;
and2_9574: n_10885 <=  n_10886  AND n_10887;
inv_9575: n_10886  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_9576: n_10887  <= TRANSPORT a_SCH0ADDRREG_F14_G  ;
and1_9577: n_10888 <=  gnd;
delay_9578: a_N240_aNOT  <= TRANSPORT a_EQ219  ;
xor2_9579: a_EQ219 <=  n_10891  XOR n_10898;
or2_9580: n_10891 <=  n_10892  OR n_10895;
and2_9581: n_10892 <=  n_10893  AND n_10894;
inv_9582: n_10893  <= TRANSPORT NOT a_N2531  ;
delay_9583: n_10894  <= TRANSPORT a_LC4_F9  ;
and2_9584: n_10895 <=  n_10896  AND n_10897;
delay_9585: n_10896  <= TRANSPORT a_N2531  ;
delay_9586: n_10897  <= TRANSPORT a_LC7_F9  ;
and1_9587: n_10898 <=  gnd;
delay_9588: a_LC3_F9  <= TRANSPORT a_EQ216  ;
xor2_9589: a_EQ216 <=  n_10901  XOR n_10908;
or2_9590: n_10901 <=  n_10902  OR n_10905;
and2_9591: n_10902 <=  n_10903  AND n_10904;
inv_9592: n_10903  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_9593: n_10904  <= TRANSPORT a_SCH0ADDRREG_F14_G  ;
and2_9594: n_10905 <=  n_10906  AND n_10907;
inv_9595: n_10906  <= TRANSPORT NOT a_N2376  ;
delay_9596: n_10907  <= TRANSPORT a_SCH2ADDRREG_F14_G  ;
and1_9597: n_10908 <=  gnd;
delay_9598: a_LC1_F9  <= TRANSPORT a_EQ215  ;
xor2_9599: a_EQ215 <=  n_10911  XOR n_10918;
or2_9600: n_10911 <=  n_10912  OR n_10915;
and2_9601: n_10912 <=  n_10913  AND n_10914;
inv_9602: n_10913  <= TRANSPORT NOT a_N88_aNOT  ;
delay_9603: n_10914  <= TRANSPORT a_SCH1ADDRREG_F14_G  ;
and2_9604: n_10915 <=  n_10916  AND n_10917;
inv_9605: n_10916  <= TRANSPORT NOT a_N2377  ;
delay_9606: n_10917  <= TRANSPORT a_SCH3ADDRREG_F14_G  ;
and1_9607: n_10918 <=  gnd;
dff_9608: DFF_a8237

    PORT MAP ( D => a_EQ860, CLK => a_SADDRESSOUT_F14_G_aCLK, CLRN => a_SADDRESSOUT_F14_G_aCLRN,
          PRN => vcc, Q => a_SADDRESSOUT_F14_G);
inv_9609: a_SADDRESSOUT_F14_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9610: a_EQ860 <=  n_10925  XOR n_10935;
or3_9611: n_10925 <=  n_10926  OR n_10929  OR n_10932;
and2_9612: n_10926 <=  n_10927  AND n_10928;
delay_9613: n_10927  <= TRANSPORT a_N240_aNOT  ;
inv_9614: n_10928  <= TRANSPORT NOT startdma  ;
and2_9615: n_10929 <=  n_10930  AND n_10931;
delay_9616: n_10930  <= TRANSPORT a_LC3_F9  ;
delay_9617: n_10931  <= TRANSPORT startdma  ;
and2_9618: n_10932 <=  n_10933  AND n_10934;
delay_9619: n_10933  <= TRANSPORT a_LC1_F9  ;
delay_9620: n_10934  <= TRANSPORT startdma  ;
and1_9621: n_10935 <=  gnd;
delay_9622: n_10936  <= TRANSPORT clk  ;
filter_9623: FILTER_a8237

    PORT MAP (IN1 => n_10936, Y => a_SADDRESSOUT_F14_G_aCLK);
delay_9624: a_N1776_aNOT  <= TRANSPORT a_EQ508  ;
xor2_9625: a_EQ508 <=  n_10940  XOR n_10947;
or2_9626: n_10940 <=  n_10941  OR n_10944;
and2_9627: n_10941 <=  n_10942  AND n_10943;
delay_9628: n_10942  <= TRANSPORT a_LC4_A3  ;
delay_9629: n_10943  <= TRANSPORT bytepointer  ;
and2_9630: n_10944 <=  n_10945  AND n_10946;
delay_9631: n_10945  <= TRANSPORT a_N87  ;
delay_9632: n_10946  <= TRANSPORT bytepointer  ;
and1_9633: n_10947 <=  gnd;
delay_9634: a_LC6_A4  <= TRANSPORT a_LC6_A4_aIN  ;
xor2_9635: a_LC6_A4_aIN <=  n_10950  XOR n_10955;
or1_9636: n_10950 <=  n_10951;
and3_9637: n_10951 <=  n_10952  AND n_10953  AND n_10954;
delay_9638: n_10952  <= TRANSPORT niowin  ;
inv_9639: n_10953  <= TRANSPORT NOT niorin  ;
inv_9640: n_10954  <= TRANSPORT NOT ncs  ;
and1_9641: n_10955 <=  gnd;
dff_9642: DFF_a8237

    PORT MAP ( D => a_EQ001, CLK => bytepointer_aCLK, CLRN => bytepointer_aCLRN,
          PRN => vcc, Q => bytepointer);
inv_9643: bytepointer_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9644: a_EQ001 <=  n_10962  XOR n_10969;
or2_9645: n_10962 <=  n_10963  OR n_10965;
and1_9646: n_10963 <=  n_10964;
delay_9647: n_10964  <= TRANSPORT a_N1776_aNOT  ;
and3_9648: n_10965 <=  n_10966  AND n_10967  AND n_10968;
inv_9649: n_10966  <= TRANSPORT NOT a_LC4_A3  ;
delay_9650: n_10967  <= TRANSPORT a_LC6_A4  ;
inv_9651: n_10968  <= TRANSPORT NOT ain(0)  ;
and1_9652: n_10969 <=  gnd;
delay_9653: n_10970  <= TRANSPORT clk  ;
filter_9654: FILTER_a8237

    PORT MAP (IN1 => n_10970, Y => bytepointer_aCLK);
dff_9655: DFF_a8237

    PORT MAP ( D => a_EQ1188, CLK => a_STEMPORARYREG_F7_G_aCLK, CLRN => a_STEMPORARYREG_F7_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F7_G);
inv_9656: a_STEMPORARYREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9657: a_EQ1188 <=  n_10979  XOR n_10988;
or2_9658: n_10979 <=  n_10980  OR n_10984;
and3_9659: n_10980 <=  n_10981  AND n_10982  AND n_10983;
delay_9660: n_10981  <= TRANSPORT a_N2563_aNOT  ;
inv_9661: n_10982  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_9662: n_10983  <= TRANSPORT a_STEMPORARYREG_F7_G  ;
and3_9663: n_10984 <=  n_10985  AND n_10986  AND n_10987;
delay_9664: n_10985  <= TRANSPORT a_N2563_aNOT  ;
delay_9665: n_10986  <= TRANSPORT a_N2372_aNOT  ;
delay_9666: n_10987  <= TRANSPORT dbin(7)  ;
and1_9667: n_10988 <=  gnd;
delay_9668: n_10989  <= TRANSPORT clk  ;
filter_9669: FILTER_a8237

    PORT MAP (IN1 => n_10989, Y => a_STEMPORARYREG_F7_G_aCLK);
delay_9670: a_LC2_F19  <= TRANSPORT a_EQ285  ;
xor2_9671: a_EQ285 <=  n_10993  XOR n_11005;
or3_9672: n_10993 <=  n_10994  OR n_10998  OR n_11001;
and2_9673: n_10994 <=  n_10995  AND n_10996;
delay_9674: n_10995  <= TRANSPORT a_N77_aNOT  ;
delay_9675: n_10996  <= TRANSPORT a_SCH2ADDRREG_F0_G  ;
and2_9676: n_10998 <=  n_10999  AND n_11000;
delay_9677: n_10999  <= TRANSPORT a_LC6_D6  ;
delay_9678: n_11000  <= TRANSPORT a_SCH2ADDRREG_F0_G  ;
and3_9679: n_11001 <=  n_11002  AND n_11003  AND n_11004;
inv_9680: n_11002  <= TRANSPORT NOT a_LC6_D6  ;
inv_9681: n_11003  <= TRANSPORT NOT a_N77_aNOT  ;
delay_9682: n_11004  <= TRANSPORT dbin(0)  ;
and1_9683: n_11005 <=  gnd;
delay_9684: a_LC3_F19  <= TRANSPORT a_EQ723  ;
xor2_9685: a_EQ723 <=  n_11008  XOR n_11019;
or3_9686: n_11008 <=  n_11009  OR n_11013  OR n_11016;
and3_9687: n_11009 <=  n_11010  AND n_11011  AND n_11012;
delay_9688: n_11010  <= TRANSPORT a_N2557  ;
inv_9689: n_11011  <= TRANSPORT NOT a_N2376  ;
inv_9690: n_11012  <= TRANSPORT NOT a_LC7_D18  ;
and2_9691: n_11013 <=  n_11014  AND n_11015;
inv_9692: n_11014  <= TRANSPORT NOT a_N2557  ;
delay_9693: n_11015  <= TRANSPORT a_LC2_F19  ;
and2_9694: n_11016 <=  n_11017  AND n_11018;
delay_9695: n_11017  <= TRANSPORT a_N2376  ;
delay_9696: n_11018  <= TRANSPORT a_LC2_F19  ;
and1_9697: n_11019 <=  gnd;
dff_9698: DFF_a8237

    PORT MAP ( D => a_EQ995, CLK => a_SCH2ADDRREG_F0_G_aCLK, CLRN => a_SCH2ADDRREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F0_G);
inv_9699: a_SCH2ADDRREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9700: a_EQ995 <=  n_11026  XOR n_11037;
or3_9701: n_11026 <=  n_11027  OR n_11031  OR n_11034;
and3_9702: n_11027 <=  n_11028  AND n_11029  AND n_11030;
delay_9703: n_11028  <= TRANSPORT a_N57_aNOT  ;
delay_9704: n_11029  <= TRANSPORT a_SCH2BAROUT_F0_G  ;
delay_9705: n_11030  <= TRANSPORT a_SCH2MODEREG_F2_G  ;
and2_9706: n_11031 <=  n_11032  AND n_11033;
inv_9707: n_11032  <= TRANSPORT NOT a_SCH2MODEREG_F2_G  ;
delay_9708: n_11033  <= TRANSPORT a_LC3_F19  ;
and2_9709: n_11034 <=  n_11035  AND n_11036;
inv_9710: n_11035  <= TRANSPORT NOT a_N57_aNOT  ;
delay_9711: n_11036  <= TRANSPORT a_LC3_F19  ;
and1_9712: n_11037 <=  gnd;
delay_9713: n_11038  <= TRANSPORT clk  ;
filter_9714: FILTER_a8237

    PORT MAP (IN1 => n_11038, Y => a_SCH2ADDRREG_F0_G_aCLK);
delay_9715: a_N1493_aNOT  <= TRANSPORT a_EQ455  ;
xor2_9716: a_EQ455 <=  n_11042  XOR n_11054;
or3_9717: n_11042 <=  n_11043  OR n_11047  OR n_11050;
and2_9718: n_11043 <=  n_11044  AND n_11045;
delay_9719: n_11044  <= TRANSPORT a_N2348  ;
delay_9720: n_11045  <= TRANSPORT a_SCH3ADDRREG_F0_G  ;
and2_9721: n_11047 <=  n_11048  AND n_11049;
delay_9722: n_11048  <= TRANSPORT a_LC6_D6  ;
delay_9723: n_11049  <= TRANSPORT a_SCH3ADDRREG_F0_G  ;
and3_9724: n_11050 <=  n_11051  AND n_11052  AND n_11053;
inv_9725: n_11051  <= TRANSPORT NOT a_LC6_D6  ;
inv_9726: n_11052  <= TRANSPORT NOT a_N2348  ;
delay_9727: n_11053  <= TRANSPORT dbin(0)  ;
and1_9728: n_11054 <=  gnd;
delay_9729: a_LC8_D8  <= TRANSPORT a_EQ456  ;
xor2_9730: a_EQ456 <=  n_11057  XOR n_11068;
or3_9731: n_11057 <=  n_11058  OR n_11062  OR n_11065;
and3_9732: n_11058 <=  n_11059  AND n_11060  AND n_11061;
delay_9733: n_11059  <= TRANSPORT a_N2557  ;
inv_9734: n_11060  <= TRANSPORT NOT a_N2377  ;
inv_9735: n_11061  <= TRANSPORT NOT a_LC7_D18  ;
and2_9736: n_11062 <=  n_11063  AND n_11064;
inv_9737: n_11063  <= TRANSPORT NOT a_N2557  ;
delay_9738: n_11064  <= TRANSPORT a_N1493_aNOT  ;
and2_9739: n_11065 <=  n_11066  AND n_11067;
delay_9740: n_11066  <= TRANSPORT a_N2377  ;
delay_9741: n_11067  <= TRANSPORT a_N1493_aNOT  ;
and1_9742: n_11068 <=  gnd;
dff_9743: DFF_a8237

    PORT MAP ( D => a_EQ1059, CLK => a_SCH3ADDRREG_F0_G_aCLK, CLRN => a_SCH3ADDRREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F0_G);
inv_9744: a_SCH3ADDRREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9745: a_EQ1059 <=  n_11075  XOR n_11086;
or3_9746: n_11075 <=  n_11076  OR n_11080  OR n_11083;
and3_9747: n_11076 <=  n_11077  AND n_11078  AND n_11079;
delay_9748: n_11077  <= TRANSPORT a_N57_aNOT  ;
delay_9749: n_11078  <= TRANSPORT a_SCH3BAROUT_F0_G  ;
delay_9750: n_11079  <= TRANSPORT a_SCH3MODEREG_F2_G  ;
and2_9751: n_11080 <=  n_11081  AND n_11082;
inv_9752: n_11081  <= TRANSPORT NOT a_SCH3MODEREG_F2_G  ;
delay_9753: n_11082  <= TRANSPORT a_LC8_D8  ;
and2_9754: n_11083 <=  n_11084  AND n_11085;
inv_9755: n_11084  <= TRANSPORT NOT a_N57_aNOT  ;
delay_9756: n_11085  <= TRANSPORT a_LC8_D8  ;
and1_9757: n_11086 <=  gnd;
delay_9758: n_11087  <= TRANSPORT clk  ;
filter_9759: FILTER_a8237

    PORT MAP (IN1 => n_11087, Y => a_SCH3ADDRREG_F0_G_aCLK);
delay_9760: a_LC1_D8  <= TRANSPORT a_EQ673  ;
xor2_9761: a_EQ673 <=  n_11091  XOR n_11103;
or3_9762: n_11091 <=  n_11092  OR n_11096  OR n_11099;
and2_9763: n_11092 <=  n_11093  AND n_11094;
inv_9764: n_11093  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_9765: n_11094  <= TRANSPORT a_SCH0ADDRREG_F0_G  ;
and2_9766: n_11096 <=  n_11097  AND n_11098;
delay_9767: n_11097  <= TRANSPORT a_LC6_D6  ;
delay_9768: n_11098  <= TRANSPORT a_SCH0ADDRREG_F0_G  ;
and3_9769: n_11099 <=  n_11100  AND n_11101  AND n_11102;
inv_9770: n_11100  <= TRANSPORT NOT a_LC6_D6  ;
delay_9771: n_11101  <= TRANSPORT a_N2354_aNOT  ;
delay_9772: n_11102  <= TRANSPORT dbin(0)  ;
and1_9773: n_11103 <=  gnd;
delay_9774: a_LC4_D8  <= TRANSPORT a_EQ674  ;
xor2_9775: a_EQ674 <=  n_11106  XOR n_11118;
or3_9776: n_11106 <=  n_11107  OR n_11111  OR n_11115;
and3_9777: n_11107 <=  n_11108  AND n_11109  AND n_11110;
inv_9778: n_11108  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_9779: n_11109  <= TRANSPORT a_N2530_aNOT  ;
inv_9780: n_11110  <= TRANSPORT NOT a_LC7_D18  ;
and3_9781: n_11111 <=  n_11112  AND n_11113  AND n_11114;
inv_9782: n_11112  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_9783: n_11113  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_9784: n_11114  <= TRANSPORT a_LC7_D18  ;
and2_9785: n_11115 <=  n_11116  AND n_11117;
delay_9786: n_11116  <= TRANSPORT a_N2558_aNOT  ;
delay_9787: n_11117  <= TRANSPORT a_LC1_D8  ;
and1_9788: n_11118 <=  gnd;
dff_9789: DFF_a8237

    PORT MAP ( D => a_EQ867, CLK => a_SCH0ADDRREG_F0_G_aCLK, CLRN => a_SCH0ADDRREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F0_G);
inv_9790: a_SCH0ADDRREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9791: a_EQ867 <=  n_11125  XOR n_11136;
or3_9792: n_11125 <=  n_11126  OR n_11130  OR n_11133;
and3_9793: n_11126 <=  n_11127  AND n_11128  AND n_11129;
delay_9794: n_11127  <= TRANSPORT a_N57_aNOT  ;
delay_9795: n_11128  <= TRANSPORT a_SCH0BAROUT_F0_G  ;
delay_9796: n_11129  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and2_9797: n_11130 <=  n_11131  AND n_11132;
inv_9798: n_11131  <= TRANSPORT NOT a_SCH0MODEREG_F2_G  ;
delay_9799: n_11132  <= TRANSPORT a_LC4_D8  ;
and2_9800: n_11133 <=  n_11134  AND n_11135;
inv_9801: n_11134  <= TRANSPORT NOT a_N57_aNOT  ;
delay_9802: n_11135  <= TRANSPORT a_LC4_D8  ;
and1_9803: n_11136 <=  gnd;
delay_9804: n_11137  <= TRANSPORT clk  ;
filter_9805: FILTER_a8237

    PORT MAP (IN1 => n_11137, Y => a_SCH0ADDRREG_F0_G_aCLK);
delay_9806: a_LC2_D19  <= TRANSPORT a_EQ698  ;
xor2_9807: a_EQ698 <=  n_11141  XOR n_11153;
or3_9808: n_11141 <=  n_11142  OR n_11146  OR n_11149;
and2_9809: n_11142 <=  n_11143  AND n_11144;
delay_9810: n_11143  <= TRANSPORT a_N2352  ;
delay_9811: n_11144  <= TRANSPORT a_SCH1ADDRREG_F0_G  ;
and2_9812: n_11146 <=  n_11147  AND n_11148;
delay_9813: n_11147  <= TRANSPORT a_LC6_D6  ;
delay_9814: n_11148  <= TRANSPORT a_SCH1ADDRREG_F0_G  ;
and3_9815: n_11149 <=  n_11150  AND n_11151  AND n_11152;
inv_9816: n_11150  <= TRANSPORT NOT a_LC6_D6  ;
inv_9817: n_11151  <= TRANSPORT NOT a_N2352  ;
delay_9818: n_11152  <= TRANSPORT dbin(0)  ;
and1_9819: n_11153 <=  gnd;
delay_9820: a_LC1_D19  <= TRANSPORT a_EQ699  ;
xor2_9821: a_EQ699 <=  n_11156  XOR n_11168;
or3_9822: n_11156 <=  n_11157  OR n_11161  OR n_11165;
and3_9823: n_11157 <=  n_11158  AND n_11159  AND n_11160;
inv_9824: n_11158  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_9825: n_11159  <= TRANSPORT a_N2530_aNOT  ;
inv_9826: n_11160  <= TRANSPORT NOT a_LC7_D18  ;
and3_9827: n_11161 <=  n_11162  AND n_11163  AND n_11164;
inv_9828: n_11162  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_9829: n_11163  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_9830: n_11164  <= TRANSPORT a_LC7_D18  ;
and2_9831: n_11165 <=  n_11166  AND n_11167;
delay_9832: n_11166  <= TRANSPORT a_N2559_aNOT  ;
delay_9833: n_11167  <= TRANSPORT a_LC2_D19  ;
and1_9834: n_11168 <=  gnd;
dff_9835: DFF_a8237

    PORT MAP ( D => a_EQ931, CLK => a_SCH1ADDRREG_F0_G_aCLK, CLRN => a_SCH1ADDRREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F0_G);
inv_9836: a_SCH1ADDRREG_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9837: a_EQ931 <=  n_11175  XOR n_11186;
or3_9838: n_11175 <=  n_11176  OR n_11180  OR n_11183;
and3_9839: n_11176 <=  n_11177  AND n_11178  AND n_11179;
delay_9840: n_11177  <= TRANSPORT a_N57_aNOT  ;
delay_9841: n_11178  <= TRANSPORT a_SCH1BAROUT_F0_G  ;
delay_9842: n_11179  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and2_9843: n_11180 <=  n_11181  AND n_11182;
inv_9844: n_11181  <= TRANSPORT NOT a_SCH1MODEREG_F2_G  ;
delay_9845: n_11182  <= TRANSPORT a_LC1_D19  ;
and2_9846: n_11183 <=  n_11184  AND n_11185;
inv_9847: n_11184  <= TRANSPORT NOT a_N57_aNOT  ;
delay_9848: n_11185  <= TRANSPORT a_LC1_D19  ;
and1_9849: n_11186 <=  gnd;
delay_9850: n_11187  <= TRANSPORT clk  ;
filter_9851: FILTER_a8237

    PORT MAP (IN1 => n_11187, Y => a_SCH1ADDRREG_F0_G_aCLK);
delay_9852: a_N3059  <= TRANSPORT a_EQ836  ;
xor2_9853: a_EQ836 <=  n_11191  XOR n_11208;
or4_9854: n_11191 <=  n_11192  OR n_11196  OR n_11200  OR n_11204;
and3_9855: n_11192 <=  n_11193  AND n_11194  AND n_11195;
delay_9856: n_11193  <= TRANSPORT a_N2529  ;
inv_9857: n_11194  <= TRANSPORT NOT a_LC7_D18  ;
inv_9858: n_11195  <= TRANSPORT NOT a_LC7_C17  ;
and3_9859: n_11196 <=  n_11197  AND n_11198  AND n_11199;
delay_9860: n_11197  <= TRANSPORT a_N2529  ;
delay_9861: n_11198  <= TRANSPORT a_LC7_D18  ;
delay_9862: n_11199  <= TRANSPORT a_LC7_C17  ;
and3_9863: n_11200 <=  n_11201  AND n_11202  AND n_11203;
inv_9864: n_11201  <= TRANSPORT NOT a_N2529  ;
delay_9865: n_11202  <= TRANSPORT a_LC7_D18  ;
inv_9866: n_11203  <= TRANSPORT NOT a_LC7_C17  ;
and3_9867: n_11204 <=  n_11205  AND n_11206  AND n_11207;
inv_9868: n_11205  <= TRANSPORT NOT a_N2529  ;
inv_9869: n_11206  <= TRANSPORT NOT a_LC7_D18  ;
delay_9870: n_11207  <= TRANSPORT a_LC7_C17  ;
and1_9871: n_11208 <=  gnd;
delay_9872: a_LC3_C9  <= TRANSPORT a_EQ235  ;
xor2_9873: a_EQ235 <=  n_11211  XOR n_11220;
or2_9874: n_11211 <=  n_11212  OR n_11216;
and3_9875: n_11212 <=  n_11213  AND n_11214  AND n_11215;
inv_9876: n_11213  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_9877: n_11214  <= TRANSPORT a_N2530_aNOT  ;
delay_9878: n_11215  <= TRANSPORT a_N3059  ;
and3_9879: n_11216 <=  n_11217  AND n_11218  AND n_11219;
inv_9880: n_11217  <= TRANSPORT NOT a_N2559_aNOT  ;
inv_9881: n_11218  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_9882: n_11219  <= TRANSPORT a_LC7_C17  ;
and1_9883: n_11220 <=  gnd;
delay_9884: a_LC2_C9  <= TRANSPORT a_EQ697  ;
xor2_9885: a_EQ697 <=  n_11223  XOR n_11233;
or2_9886: n_11223 <=  n_11224  OR n_11228;
and3_9887: n_11224 <=  n_11225  AND n_11226  AND n_11227;
delay_9888: n_11225  <= TRANSPORT a_N2559_aNOT  ;
delay_9889: n_11226  <= TRANSPORT dbin(1)  ;
inv_9890: n_11227  <= TRANSPORT NOT a_N2584_aNOT  ;
and3_9891: n_11228 <=  n_11229  AND n_11230  AND n_11231;
delay_9892: n_11229  <= TRANSPORT a_N2559_aNOT  ;
delay_9893: n_11230  <= TRANSPORT a_N2584_aNOT  ;
delay_9894: n_11231  <= TRANSPORT a_SCH1ADDRREG_F1_G  ;
and1_9895: n_11233 <=  gnd;
dff_9896: DFF_a8237

    PORT MAP ( D => a_EQ932, CLK => a_SCH1ADDRREG_F1_G_aCLK, CLRN => a_SCH1ADDRREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F1_G);
inv_9897: a_SCH1ADDRREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9898: a_EQ932 <=  n_11240  XOR n_11250;
or3_9899: n_11240 <=  n_11241  OR n_11244  OR n_11247;
and2_9900: n_11241 <=  n_11242  AND n_11243;
delay_9901: n_11242  <= TRANSPORT a_N2526  ;
delay_9902: n_11243  <= TRANSPORT a_SCH1BAROUT_F1_G  ;
and2_9903: n_11244 <=  n_11245  AND n_11246;
inv_9904: n_11245  <= TRANSPORT NOT a_N2526  ;
delay_9905: n_11246  <= TRANSPORT a_LC3_C9  ;
and2_9906: n_11247 <=  n_11248  AND n_11249;
inv_9907: n_11248  <= TRANSPORT NOT a_N2526  ;
delay_9908: n_11249  <= TRANSPORT a_LC2_C9  ;
and1_9909: n_11250 <=  gnd;
delay_9910: n_11251  <= TRANSPORT clk  ;
filter_9911: FILTER_a8237

    PORT MAP (IN1 => n_11251, Y => a_SCH1ADDRREG_F1_G_aCLK);
delay_9912: a_LC4_C9  <= TRANSPORT a_EQ270  ;
xor2_9913: a_EQ270 <=  n_11255  XOR n_11264;
or2_9914: n_11255 <=  n_11256  OR n_11260;
and3_9915: n_11256 <=  n_11257  AND n_11258  AND n_11259;
inv_9916: n_11257  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_9917: n_11258  <= TRANSPORT a_N2530_aNOT  ;
delay_9918: n_11259  <= TRANSPORT a_N3059  ;
and3_9919: n_11260 <=  n_11261  AND n_11262  AND n_11263;
inv_9920: n_11261  <= TRANSPORT NOT a_N2558_aNOT  ;
inv_9921: n_11262  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_9922: n_11263  <= TRANSPORT a_LC7_C17  ;
and1_9923: n_11264 <=  gnd;
delay_9924: a_LC5_C9  <= TRANSPORT a_EQ672  ;
xor2_9925: a_EQ672 <=  n_11267  XOR n_11277;
or2_9926: n_11267 <=  n_11268  OR n_11272;
and3_9927: n_11268 <=  n_11269  AND n_11270  AND n_11271;
delay_9928: n_11269  <= TRANSPORT a_N2586  ;
delay_9929: n_11270  <= TRANSPORT a_N2558_aNOT  ;
delay_9930: n_11271  <= TRANSPORT dbin(1)  ;
and3_9931: n_11272 <=  n_11273  AND n_11274  AND n_11275;
inv_9932: n_11273  <= TRANSPORT NOT a_N2586  ;
delay_9933: n_11274  <= TRANSPORT a_N2558_aNOT  ;
delay_9934: n_11275  <= TRANSPORT a_SCH0ADDRREG_F1_G  ;
and1_9935: n_11277 <=  gnd;
dff_9936: DFF_a8237

    PORT MAP ( D => a_EQ868, CLK => a_SCH0ADDRREG_F1_G_aCLK, CLRN => a_SCH0ADDRREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F1_G);
inv_9937: a_SCH0ADDRREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9938: a_EQ868 <=  n_11284  XOR n_11294;
or3_9939: n_11284 <=  n_11285  OR n_11288  OR n_11291;
and2_9940: n_11285 <=  n_11286  AND n_11287;
delay_9941: n_11286  <= TRANSPORT a_N2525  ;
delay_9942: n_11287  <= TRANSPORT a_SCH0BAROUT_F1_G  ;
and2_9943: n_11288 <=  n_11289  AND n_11290;
inv_9944: n_11289  <= TRANSPORT NOT a_N2525  ;
delay_9945: n_11290  <= TRANSPORT a_LC4_C9  ;
and2_9946: n_11291 <=  n_11292  AND n_11293;
inv_9947: n_11292  <= TRANSPORT NOT a_N2525  ;
delay_9948: n_11293  <= TRANSPORT a_LC5_C9  ;
and1_9949: n_11294 <=  gnd;
delay_9950: n_11295  <= TRANSPORT clk  ;
filter_9951: FILTER_a8237

    PORT MAP (IN1 => n_11295, Y => a_SCH0ADDRREG_F1_G_aCLK);
delay_9952: a_LC3_C12  <= TRANSPORT a_EQ721  ;
xor2_9953: a_EQ721 <=  n_11299  XOR n_11307;
or2_9954: n_11299 <=  n_11300  OR n_11303;
and2_9955: n_11300 <=  n_11301  AND n_11302;
inv_9956: n_11301  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_9957: n_11302  <= TRANSPORT a_N3059  ;
and3_9958: n_11303 <=  n_11304  AND n_11305  AND n_11306;
delay_9959: n_11304  <= TRANSPORT a_N2560_aNOT  ;
inv_9960: n_11305  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_9961: n_11306  <= TRANSPORT dbin(1)  ;
and1_9962: n_11307 <=  gnd;
delay_9963: a_LC5_C12  <= TRANSPORT a_EQ722  ;
xor2_9964: a_EQ722 <=  n_11310  XOR n_11317;
or2_9965: n_11310 <=  n_11311  OR n_11314;
and2_9966: n_11311 <=  n_11312  AND n_11313;
delay_9967: n_11312  <= TRANSPORT a_N2527  ;
delay_9968: n_11313  <= TRANSPORT a_SCH2BAROUT_F1_G  ;
and2_9969: n_11314 <=  n_11315  AND n_11316;
inv_9970: n_11315  <= TRANSPORT NOT a_N2527  ;
delay_9971: n_11316  <= TRANSPORT a_LC3_C12  ;
and1_9972: n_11317 <=  gnd;
dff_9973: DFF_a8237

    PORT MAP ( D => a_EQ996, CLK => a_SCH2ADDRREG_F1_G_aCLK, CLRN => a_SCH2ADDRREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F1_G);
inv_9974: a_SCH2ADDRREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_9975: a_EQ996 <=  n_11325  XOR n_11332;
or2_9976: n_11325 <=  n_11326  OR n_11328;
and1_9977: n_11326 <=  n_11327;
delay_9978: n_11327  <= TRANSPORT a_LC5_C12  ;
and3_9979: n_11328 <=  n_11329  AND n_11330  AND n_11331;
delay_9980: n_11329  <= TRANSPORT a_N756  ;
delay_9981: n_11330  <= TRANSPORT a_N2582_aNOT  ;
delay_9982: n_11331  <= TRANSPORT a_SCH2ADDRREG_F1_G  ;
and1_9983: n_11332 <=  gnd;
delay_9984: n_11333  <= TRANSPORT clk  ;
filter_9985: FILTER_a8237

    PORT MAP (IN1 => n_11333, Y => a_SCH2ADDRREG_F1_G_aCLK);
delay_9986: a_N937_aNOT  <= TRANSPORT a_N937_aNOT_aIN  ;
xor2_9987: a_N937_aNOT_aIN <=  n_11337  XOR n_11341;
or1_9988: n_11337 <=  n_11338;
and2_9989: n_11338 <=  n_11339  AND n_11340;
delay_9990: n_11339  <= TRANSPORT a_N1094  ;
delay_9991: n_11340  <= TRANSPORT a_N3059  ;
and1_9992: n_11341 <=  gnd;
delay_9993: a_LC2_C26  <= TRANSPORT a_EQ747  ;
xor2_9994: a_EQ747 <=  n_11344  XOR n_11354;
or2_9995: n_11344 <=  n_11345  OR n_11349;
and3_9996: n_11345 <=  n_11346  AND n_11347  AND n_11348;
delay_9997: n_11346  <= TRANSPORT a_N1095  ;
inv_9998: n_11347  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_9999: n_11348  <= TRANSPORT dbin(1)  ;
and3_10000: n_11349 <=  n_11350  AND n_11351  AND n_11352;
delay_10001: n_11350  <= TRANSPORT a_N1095  ;
delay_10002: n_11351  <= TRANSPORT a_N2580_aNOT  ;
delay_10003: n_11352  <= TRANSPORT a_SCH3ADDRREG_F1_G  ;
and1_10004: n_11354 <=  gnd;
dff_10005: DFF_a8237

    PORT MAP ( D => a_EQ1060, CLK => a_SCH3ADDRREG_F1_G_aCLK, CLRN => a_SCH3ADDRREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F1_G);
inv_10006: a_SCH3ADDRREG_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10007: a_EQ1060 <=  n_11361  XOR n_11369;
or3_10008: n_11361 <=  n_11362  OR n_11364  OR n_11366;
and1_10009: n_11362 <=  n_11363;
delay_10010: n_11363  <= TRANSPORT a_N937_aNOT  ;
and1_10011: n_11364 <=  n_11365;
delay_10012: n_11365  <= TRANSPORT a_LC2_C26  ;
and2_10013: n_11366 <=  n_11367  AND n_11368;
delay_10014: n_11367  <= TRANSPORT a_N2528  ;
delay_10015: n_11368  <= TRANSPORT a_SCH3BAROUT_F1_G  ;
and1_10016: n_11369 <=  gnd;
delay_10017: n_11370  <= TRANSPORT clk  ;
filter_10018: FILTER_a8237

    PORT MAP (IN1 => n_11370, Y => a_SCH3ADDRREG_F1_G_aCLK);
delay_10019: a_N2542  <= TRANSPORT a_EQ599  ;
xor2_10020: a_EQ599 <=  n_11374  XOR n_11386;
or3_10021: n_11374 <=  n_11375  OR n_11379  OR n_11383;
and3_10022: n_11375 <=  n_11376  AND n_11377  AND n_11378;
inv_10023: n_11376  <= TRANSPORT NOT a_N2529  ;
delay_10024: n_11377  <= TRANSPORT a_N2530_aNOT  ;
delay_10025: n_11378  <= TRANSPORT a_LC2_C14  ;
and3_10026: n_11379 <=  n_11380  AND n_11381  AND n_11382;
delay_10027: n_11380  <= TRANSPORT a_N2529  ;
delay_10028: n_11381  <= TRANSPORT a_N2530_aNOT  ;
inv_10029: n_11382  <= TRANSPORT NOT a_LC2_C14  ;
and2_10030: n_11383 <=  n_11384  AND n_11385;
inv_10031: n_11384  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_10032: n_11385  <= TRANSPORT a_LC4_C16  ;
and1_10033: n_11386 <=  gnd;
delay_10034: a_LC1_C2  <= TRANSPORT a_EQ695  ;
xor2_10035: a_EQ695 <=  n_11389  XOR n_11401;
or3_10036: n_11389 <=  n_11390  OR n_11394  OR n_11397;
and2_10037: n_11390 <=  n_11391  AND n_11392;
delay_10038: n_11391  <= TRANSPORT a_N2352  ;
delay_10039: n_11392  <= TRANSPORT a_SCH1ADDRREG_F2_G  ;
and2_10040: n_11394 <=  n_11395  AND n_11396;
delay_10041: n_11395  <= TRANSPORT a_LC6_D6  ;
delay_10042: n_11396  <= TRANSPORT a_SCH1ADDRREG_F2_G  ;
and3_10043: n_11397 <=  n_11398  AND n_11399  AND n_11400;
inv_10044: n_11398  <= TRANSPORT NOT a_LC6_D6  ;
inv_10045: n_11399  <= TRANSPORT NOT a_N2352  ;
delay_10046: n_11400  <= TRANSPORT dbin(2)  ;
and1_10047: n_11401 <=  gnd;
delay_10048: a_LC2_C2  <= TRANSPORT a_EQ696  ;
xor2_10049: a_EQ696 <=  n_11404  XOR n_11411;
or2_10050: n_11404 <=  n_11405  OR n_11408;
and2_10051: n_11405 <=  n_11406  AND n_11407;
inv_10052: n_11406  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_10053: n_11407  <= TRANSPORT a_N2542  ;
and2_10054: n_11408 <=  n_11409  AND n_11410;
delay_10055: n_11409  <= TRANSPORT a_N2559_aNOT  ;
delay_10056: n_11410  <= TRANSPORT a_LC1_C2  ;
and1_10057: n_11411 <=  gnd;
dff_10058: DFF_a8237

    PORT MAP ( D => a_EQ933, CLK => a_SCH1ADDRREG_F2_G_aCLK, CLRN => a_SCH1ADDRREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F2_G);
inv_10059: a_SCH1ADDRREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10060: a_EQ933 <=  n_11418  XOR n_11429;
or3_10061: n_11418 <=  n_11419  OR n_11422  OR n_11425;
and2_10062: n_11419 <=  n_11420  AND n_11421;
inv_10063: n_11420  <= TRANSPORT NOT a_SCH1MODEREG_F2_G  ;
delay_10064: n_11421  <= TRANSPORT a_LC2_C2  ;
and2_10065: n_11422 <=  n_11423  AND n_11424;
inv_10066: n_11423  <= TRANSPORT NOT a_N57_aNOT  ;
delay_10067: n_11424  <= TRANSPORT a_LC2_C2  ;
and3_10068: n_11425 <=  n_11426  AND n_11427  AND n_11428;
delay_10069: n_11426  <= TRANSPORT a_N57_aNOT  ;
delay_10070: n_11427  <= TRANSPORT a_SCH1BAROUT_F2_G  ;
delay_10071: n_11428  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and1_10072: n_11429 <=  gnd;
delay_10073: n_11430  <= TRANSPORT clk  ;
filter_10074: FILTER_a8237

    PORT MAP (IN1 => n_11430, Y => a_SCH1ADDRREG_F2_G_aCLK);
delay_10075: a_N930_aNOT  <= TRANSPORT a_EQ325  ;
xor2_10076: a_EQ325 <=  n_11434  XOR n_11443;
or2_10077: n_11434 <=  n_11435  OR n_11439;
and3_10078: n_11435 <=  n_11436  AND n_11437  AND n_11438;
delay_10079: n_11436  <= TRANSPORT a_N1094  ;
inv_10080: n_11437  <= TRANSPORT NOT a_N2529  ;
delay_10081: n_11438  <= TRANSPORT a_LC2_C14  ;
and3_10082: n_11439 <=  n_11440  AND n_11441  AND n_11442;
delay_10083: n_11440  <= TRANSPORT a_N1094  ;
delay_10084: n_11441  <= TRANSPORT a_N2529  ;
inv_10085: n_11442  <= TRANSPORT NOT a_LC2_C14  ;
and1_10086: n_11443 <=  gnd;
delay_10087: a_LC5_C20  <= TRANSPORT a_EQ746  ;
xor2_10088: a_EQ746 <=  n_11446  XOR n_11456;
or2_10089: n_11446 <=  n_11447  OR n_11451;
and3_10090: n_11447 <=  n_11448  AND n_11449  AND n_11450;
delay_10091: n_11448  <= TRANSPORT a_N1095  ;
inv_10092: n_11449  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_10093: n_11450  <= TRANSPORT dbin(2)  ;
and3_10094: n_11451 <=  n_11452  AND n_11453  AND n_11454;
delay_10095: n_11452  <= TRANSPORT a_N1095  ;
delay_10096: n_11453  <= TRANSPORT a_N2580_aNOT  ;
delay_10097: n_11454  <= TRANSPORT a_SCH3ADDRREG_F2_G  ;
and1_10098: n_11456 <=  gnd;
dff_10099: DFF_a8237

    PORT MAP ( D => a_EQ1061, CLK => a_SCH3ADDRREG_F2_G_aCLK, CLRN => a_SCH3ADDRREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F2_G);
inv_10100: a_SCH3ADDRREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10101: a_EQ1061 <=  n_11463  XOR n_11471;
or3_10102: n_11463 <=  n_11464  OR n_11466  OR n_11468;
and1_10103: n_11464 <=  n_11465;
delay_10104: n_11465  <= TRANSPORT a_N930_aNOT  ;
and1_10105: n_11466 <=  n_11467;
delay_10106: n_11467  <= TRANSPORT a_LC5_C20  ;
and2_10107: n_11468 <=  n_11469  AND n_11470;
delay_10108: n_11469  <= TRANSPORT a_N2528  ;
delay_10109: n_11470  <= TRANSPORT a_SCH3BAROUT_F2_G  ;
and1_10110: n_11471 <=  gnd;
delay_10111: n_11472  <= TRANSPORT clk  ;
filter_10112: FILTER_a8237

    PORT MAP (IN1 => n_11472, Y => a_SCH3ADDRREG_F2_G_aCLK);
delay_10113: a_N740_aNOT  <= TRANSPORT a_N740_aNOT_aIN  ;
xor2_10114: a_N740_aNOT_aIN <=  n_11476  XOR n_11483;
or1_10115: n_11476 <=  n_11477;
and4_10116: n_11477 <=  n_11478  AND n_11479  AND n_11480  AND n_11481;
delay_10117: n_11478  <= TRANSPORT a_N2560_aNOT  ;
inv_10118: n_11479  <= TRANSPORT NOT a_N2527  ;
delay_10119: n_11480  <= TRANSPORT a_N2582_aNOT  ;
delay_10120: n_11481  <= TRANSPORT a_SCH2ADDRREG_F2_G  ;
and1_10121: n_11483 <=  gnd;
delay_10122: a_N2434  <= TRANSPORT a_N2434_aIN  ;
xor2_10123: a_N2434_aIN <=  n_11486  XOR n_11490;
or1_10124: n_11486 <=  n_11487;
and2_10125: n_11487 <=  n_11488  AND n_11489;
inv_10126: n_11488  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_10127: n_11489  <= TRANSPORT dbin(2)  ;
and1_10128: n_11490 <=  gnd;
delay_10129: a_LC4_C5  <= TRANSPORT a_EQ720  ;
xor2_10130: a_EQ720 <=  n_11493  XOR n_11505;
or3_10131: n_11493 <=  n_11494  OR n_11498  OR n_11502;
and3_10132: n_11494 <=  n_11495  AND n_11496  AND n_11497;
inv_10133: n_11495  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10134: n_11496  <= TRANSPORT NOT a_N2529  ;
delay_10135: n_11497  <= TRANSPORT a_LC2_C14  ;
and3_10136: n_11498 <=  n_11499  AND n_11500  AND n_11501;
inv_10137: n_11499  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10138: n_11500  <= TRANSPORT a_N2529  ;
inv_10139: n_11501  <= TRANSPORT NOT a_LC2_C14  ;
and2_10140: n_11502 <=  n_11503  AND n_11504;
delay_10141: n_11503  <= TRANSPORT a_N2560_aNOT  ;
delay_10142: n_11504  <= TRANSPORT a_N2434  ;
and1_10143: n_11505 <=  gnd;
dff_10144: DFF_a8237

    PORT MAP ( D => a_EQ997, CLK => a_SCH2ADDRREG_F2_G_aCLK, CLRN => a_SCH2ADDRREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F2_G);
inv_10145: a_SCH2ADDRREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10146: a_EQ997 <=  n_11512  XOR n_11521;
or3_10147: n_11512 <=  n_11513  OR n_11515  OR n_11518;
and1_10148: n_11513 <=  n_11514;
delay_10149: n_11514  <= TRANSPORT a_N740_aNOT  ;
and2_10150: n_11515 <=  n_11516  AND n_11517;
inv_10151: n_11516  <= TRANSPORT NOT a_N2527  ;
delay_10152: n_11517  <= TRANSPORT a_LC4_C5  ;
and2_10153: n_11518 <=  n_11519  AND n_11520;
delay_10154: n_11519  <= TRANSPORT a_N2527  ;
delay_10155: n_11520  <= TRANSPORT a_SCH2BAROUT_F2_G  ;
and1_10156: n_11521 <=  gnd;
delay_10157: n_11522  <= TRANSPORT clk  ;
filter_10158: FILTER_a8237

    PORT MAP (IN1 => n_11522, Y => a_SCH2ADDRREG_F2_G_aCLK);
delay_10159: a_LC3_C2  <= TRANSPORT a_EQ670  ;
xor2_10160: a_EQ670 <=  n_11526  XOR n_11538;
or3_10161: n_11526 <=  n_11527  OR n_11531  OR n_11534;
and2_10162: n_11527 <=  n_11528  AND n_11529;
inv_10163: n_11528  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_10164: n_11529  <= TRANSPORT a_SCH0ADDRREG_F2_G  ;
and2_10165: n_11531 <=  n_11532  AND n_11533;
delay_10166: n_11532  <= TRANSPORT a_LC6_D6  ;
delay_10167: n_11533  <= TRANSPORT a_SCH0ADDRREG_F2_G  ;
and3_10168: n_11534 <=  n_11535  AND n_11536  AND n_11537;
inv_10169: n_11535  <= TRANSPORT NOT a_LC6_D6  ;
delay_10170: n_11536  <= TRANSPORT a_N2354_aNOT  ;
delay_10171: n_11537  <= TRANSPORT dbin(2)  ;
and1_10172: n_11538 <=  gnd;
delay_10173: a_LC4_C2  <= TRANSPORT a_EQ671  ;
xor2_10174: a_EQ671 <=  n_11541  XOR n_11548;
or2_10175: n_11541 <=  n_11542  OR n_11545;
and2_10176: n_11542 <=  n_11543  AND n_11544;
inv_10177: n_11543  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_10178: n_11544  <= TRANSPORT a_N2542  ;
and2_10179: n_11545 <=  n_11546  AND n_11547;
delay_10180: n_11546  <= TRANSPORT a_N2558_aNOT  ;
delay_10181: n_11547  <= TRANSPORT a_LC3_C2  ;
and1_10182: n_11548 <=  gnd;
dff_10183: DFF_a8237

    PORT MAP ( D => a_EQ869, CLK => a_SCH0ADDRREG_F2_G_aCLK, CLRN => a_SCH0ADDRREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F2_G);
inv_10184: a_SCH0ADDRREG_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10185: a_EQ869 <=  n_11555  XOR n_11566;
or3_10186: n_11555 <=  n_11556  OR n_11559  OR n_11562;
and2_10187: n_11556 <=  n_11557  AND n_11558;
inv_10188: n_11557  <= TRANSPORT NOT a_SCH0MODEREG_F2_G  ;
delay_10189: n_11558  <= TRANSPORT a_LC4_C2  ;
and2_10190: n_11559 <=  n_11560  AND n_11561;
inv_10191: n_11560  <= TRANSPORT NOT a_N57_aNOT  ;
delay_10192: n_11561  <= TRANSPORT a_LC4_C2  ;
and3_10193: n_11562 <=  n_11563  AND n_11564  AND n_11565;
delay_10194: n_11563  <= TRANSPORT a_N57_aNOT  ;
delay_10195: n_11564  <= TRANSPORT a_SCH0BAROUT_F2_G  ;
delay_10196: n_11565  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and1_10197: n_11566 <=  gnd;
delay_10198: n_11567  <= TRANSPORT clk  ;
filter_10199: FILTER_a8237

    PORT MAP (IN1 => n_11567, Y => a_SCH0ADDRREG_F2_G_aCLK);
delay_10200: a_N2543  <= TRANSPORT a_EQ600  ;
xor2_10201: a_EQ600 <=  n_11571  XOR n_11593;
or5_10202: n_11571 <=  n_11572  OR n_11576  OR n_11580  OR n_11583  OR n_11588;
and3_10203: n_11572 <=  n_11573  AND n_11574  AND n_11575;
delay_10204: n_11573  <= TRANSPORT a_N2529  ;
delay_10205: n_11574  <= TRANSPORT a_LC4_C14  ;
delay_10206: n_11575  <= TRANSPORT a_LC2_C24  ;
and3_10207: n_11576 <=  n_11577  AND n_11578  AND n_11579;
inv_10208: n_11577  <= TRANSPORT NOT a_N2529  ;
inv_10209: n_11578  <= TRANSPORT NOT a_LC4_C14  ;
delay_10210: n_11579  <= TRANSPORT a_LC2_C24  ;
and2_10211: n_11580 <=  n_11581  AND n_11582;
inv_10212: n_11581  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_10213: n_11582  <= TRANSPORT a_LC2_C24  ;
and4_10214: n_11583 <=  n_11584  AND n_11585  AND n_11586  AND n_11587;
inv_10215: n_11584  <= TRANSPORT NOT a_N2529  ;
delay_10216: n_11585  <= TRANSPORT a_N2530_aNOT  ;
delay_10217: n_11586  <= TRANSPORT a_LC4_C14  ;
inv_10218: n_11587  <= TRANSPORT NOT a_LC2_C24  ;
and4_10219: n_11588 <=  n_11589  AND n_11590  AND n_11591  AND n_11592;
delay_10220: n_11589  <= TRANSPORT a_N2529  ;
delay_10221: n_11590  <= TRANSPORT a_N2530_aNOT  ;
inv_10222: n_11591  <= TRANSPORT NOT a_LC4_C14  ;
inv_10223: n_11592  <= TRANSPORT NOT a_LC2_C24  ;
and1_10224: n_11593 <=  gnd;
delay_10225: a_LC4_C11  <= TRANSPORT a_EQ668  ;
xor2_10226: a_EQ668 <=  n_11596  XOR n_11604;
or2_10227: n_11596 <=  n_11597  OR n_11600;
and2_10228: n_11597 <=  n_11598  AND n_11599;
delay_10229: n_11598  <= TRANSPORT a_N2586  ;
delay_10230: n_11599  <= TRANSPORT dbin(3)  ;
and2_10231: n_11600 <=  n_11601  AND n_11602;
inv_10232: n_11601  <= TRANSPORT NOT a_N2586  ;
delay_10233: n_11602  <= TRANSPORT a_SCH0ADDRREG_F3_G  ;
and1_10234: n_11604 <=  gnd;
delay_10235: a_LC2_C11  <= TRANSPORT a_EQ669  ;
xor2_10236: a_EQ669 <=  n_11607  XOR n_11614;
or2_10237: n_11607 <=  n_11608  OR n_11611;
and2_10238: n_11608 <=  n_11609  AND n_11610;
inv_10239: n_11609  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_10240: n_11610  <= TRANSPORT a_N2543  ;
and2_10241: n_11611 <=  n_11612  AND n_11613;
delay_10242: n_11612  <= TRANSPORT a_N2558_aNOT  ;
delay_10243: n_11613  <= TRANSPORT a_LC4_C11  ;
and1_10244: n_11614 <=  gnd;
dff_10245: DFF_a8237

    PORT MAP ( D => a_EQ870, CLK => a_SCH0ADDRREG_F3_G_aCLK, CLRN => a_SCH0ADDRREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F3_G);
inv_10246: a_SCH0ADDRREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10247: a_EQ870 <=  n_11621  XOR n_11628;
or2_10248: n_11621 <=  n_11622  OR n_11625;
and2_10249: n_11622 <=  n_11623  AND n_11624;
inv_10250: n_11623  <= TRANSPORT NOT a_N2525  ;
delay_10251: n_11624  <= TRANSPORT a_LC2_C11  ;
and2_10252: n_11625 <=  n_11626  AND n_11627;
delay_10253: n_11626  <= TRANSPORT a_N2525  ;
delay_10254: n_11627  <= TRANSPORT a_SCH0BAROUT_F3_G  ;
and1_10255: n_11628 <=  gnd;
delay_10256: n_11629  <= TRANSPORT clk  ;
filter_10257: FILTER_a8237

    PORT MAP (IN1 => n_11629, Y => a_SCH0ADDRREG_F3_G_aCLK);
delay_10258: a_LC3_C7  <= TRANSPORT a_EQ286  ;
xor2_10259: a_EQ286 <=  n_11633  XOR n_11654;
or4_10260: n_11633 <=  n_11634  OR n_11639  OR n_11644  OR n_11649;
and4_10261: n_11634 <=  n_11635  AND n_11636  AND n_11637  AND n_11638;
inv_10262: n_11635  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10263: n_11636  <= TRANSPORT a_N2529  ;
delay_10264: n_11637  <= TRANSPORT a_LC4_C14  ;
delay_10265: n_11638  <= TRANSPORT a_LC2_C24  ;
and4_10266: n_11639 <=  n_11640  AND n_11641  AND n_11642  AND n_11643;
inv_10267: n_11640  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10268: n_11641  <= TRANSPORT a_N2529  ;
inv_10269: n_11642  <= TRANSPORT NOT a_LC4_C14  ;
inv_10270: n_11643  <= TRANSPORT NOT a_LC2_C24  ;
and4_10271: n_11644 <=  n_11645  AND n_11646  AND n_11647  AND n_11648;
inv_10272: n_11645  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10273: n_11646  <= TRANSPORT NOT a_N2529  ;
inv_10274: n_11647  <= TRANSPORT NOT a_LC4_C14  ;
delay_10275: n_11648  <= TRANSPORT a_LC2_C24  ;
and4_10276: n_11649 <=  n_11650  AND n_11651  AND n_11652  AND n_11653;
inv_10277: n_11650  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10278: n_11651  <= TRANSPORT NOT a_N2529  ;
delay_10279: n_11652  <= TRANSPORT a_LC4_C14  ;
inv_10280: n_11653  <= TRANSPORT NOT a_LC2_C24  ;
and1_10281: n_11654 <=  gnd;
delay_10282: a_LC4_C7  <= TRANSPORT a_EQ719  ;
xor2_10283: a_EQ719 <=  n_11657  XOR n_11667;
or2_10284: n_11657 <=  n_11658  OR n_11662;
and3_10285: n_11658 <=  n_11659  AND n_11660  AND n_11661;
delay_10286: n_11659  <= TRANSPORT a_N2560_aNOT  ;
inv_10287: n_11660  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_10288: n_11661  <= TRANSPORT dbin(3)  ;
and3_10289: n_11662 <=  n_11663  AND n_11664  AND n_11665;
delay_10290: n_11663  <= TRANSPORT a_N2560_aNOT  ;
delay_10291: n_11664  <= TRANSPORT a_N2582_aNOT  ;
delay_10292: n_11665  <= TRANSPORT a_SCH2ADDRREG_F3_G  ;
and1_10293: n_11667 <=  gnd;
dff_10294: DFF_a8237

    PORT MAP ( D => a_EQ998, CLK => a_SCH2ADDRREG_F3_G_aCLK, CLRN => a_SCH2ADDRREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F3_G);
inv_10295: a_SCH2ADDRREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10296: a_EQ998 <=  n_11674  XOR n_11684;
or3_10297: n_11674 <=  n_11675  OR n_11678  OR n_11681;
and2_10298: n_11675 <=  n_11676  AND n_11677;
inv_10299: n_11676  <= TRANSPORT NOT a_N2527  ;
delay_10300: n_11677  <= TRANSPORT a_LC3_C7  ;
and2_10301: n_11678 <=  n_11679  AND n_11680;
inv_10302: n_11679  <= TRANSPORT NOT a_N2527  ;
delay_10303: n_11680  <= TRANSPORT a_LC4_C7  ;
and2_10304: n_11681 <=  n_11682  AND n_11683;
delay_10305: n_11682  <= TRANSPORT a_N2527  ;
delay_10306: n_11683  <= TRANSPORT a_SCH2BAROUT_F3_G  ;
and1_10307: n_11684 <=  gnd;
delay_10308: n_11685  <= TRANSPORT clk  ;
filter_10309: FILTER_a8237

    PORT MAP (IN1 => n_11685, Y => a_SCH2ADDRREG_F3_G_aCLK);
delay_10310: a_LC4_C23  <= TRANSPORT a_EQ693  ;
xor2_10311: a_EQ693 <=  n_11689  XOR n_11697;
or2_10312: n_11689 <=  n_11690  OR n_11693;
and2_10313: n_11690 <=  n_11691  AND n_11692;
delay_10314: n_11691  <= TRANSPORT dbin(3)  ;
inv_10315: n_11692  <= TRANSPORT NOT a_N2584_aNOT  ;
and2_10316: n_11693 <=  n_11694  AND n_11695;
delay_10317: n_11694  <= TRANSPORT a_N2584_aNOT  ;
delay_10318: n_11695  <= TRANSPORT a_SCH1ADDRREG_F3_G  ;
and1_10319: n_11697 <=  gnd;
delay_10320: a_LC5_C23  <= TRANSPORT a_EQ694  ;
xor2_10321: a_EQ694 <=  n_11700  XOR n_11707;
or2_10322: n_11700 <=  n_11701  OR n_11704;
and2_10323: n_11701 <=  n_11702  AND n_11703;
inv_10324: n_11702  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_10325: n_11703  <= TRANSPORT a_N2543  ;
and2_10326: n_11704 <=  n_11705  AND n_11706;
delay_10327: n_11705  <= TRANSPORT a_N2559_aNOT  ;
delay_10328: n_11706  <= TRANSPORT a_LC4_C23  ;
and1_10329: n_11707 <=  gnd;
dff_10330: DFF_a8237

    PORT MAP ( D => a_EQ934, CLK => a_SCH1ADDRREG_F3_G_aCLK, CLRN => a_SCH1ADDRREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F3_G);
inv_10331: a_SCH1ADDRREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10332: a_EQ934 <=  n_11714  XOR n_11721;
or2_10333: n_11714 <=  n_11715  OR n_11718;
and2_10334: n_11715 <=  n_11716  AND n_11717;
inv_10335: n_11716  <= TRANSPORT NOT a_N2526  ;
delay_10336: n_11717  <= TRANSPORT a_LC5_C23  ;
and2_10337: n_11718 <=  n_11719  AND n_11720;
delay_10338: n_11719  <= TRANSPORT a_N2526  ;
delay_10339: n_11720  <= TRANSPORT a_SCH1BAROUT_F3_G  ;
and1_10340: n_11721 <=  gnd;
delay_10341: n_11722  <= TRANSPORT clk  ;
filter_10342: FILTER_a8237

    PORT MAP (IN1 => n_11722, Y => a_SCH1ADDRREG_F3_G_aCLK);
delay_10343: a_N944_aNOT  <= TRANSPORT a_EQ329  ;
xor2_10344: a_EQ329 <=  n_11726  XOR n_11747;
or4_10345: n_11726 <=  n_11727  OR n_11732  OR n_11737  OR n_11742;
and4_10346: n_11727 <=  n_11728  AND n_11729  AND n_11730  AND n_11731;
delay_10347: n_11728  <= TRANSPORT a_N1094  ;
delay_10348: n_11729  <= TRANSPORT a_N2529  ;
delay_10349: n_11730  <= TRANSPORT a_LC4_C14  ;
delay_10350: n_11731  <= TRANSPORT a_LC2_C24  ;
and4_10351: n_11732 <=  n_11733  AND n_11734  AND n_11735  AND n_11736;
delay_10352: n_11733  <= TRANSPORT a_N1094  ;
delay_10353: n_11734  <= TRANSPORT a_N2529  ;
inv_10354: n_11735  <= TRANSPORT NOT a_LC4_C14  ;
inv_10355: n_11736  <= TRANSPORT NOT a_LC2_C24  ;
and4_10356: n_11737 <=  n_11738  AND n_11739  AND n_11740  AND n_11741;
delay_10357: n_11738  <= TRANSPORT a_N1094  ;
inv_10358: n_11739  <= TRANSPORT NOT a_N2529  ;
inv_10359: n_11740  <= TRANSPORT NOT a_LC4_C14  ;
delay_10360: n_11741  <= TRANSPORT a_LC2_C24  ;
and4_10361: n_11742 <=  n_11743  AND n_11744  AND n_11745  AND n_11746;
delay_10362: n_11743  <= TRANSPORT a_N1094  ;
inv_10363: n_11744  <= TRANSPORT NOT a_N2529  ;
delay_10364: n_11745  <= TRANSPORT a_LC4_C14  ;
inv_10365: n_11746  <= TRANSPORT NOT a_LC2_C24  ;
and1_10366: n_11747 <=  gnd;
delay_10367: a_LC3_C26  <= TRANSPORT a_EQ745  ;
xor2_10368: a_EQ745 <=  n_11750  XOR n_11760;
or2_10369: n_11750 <=  n_11751  OR n_11755;
and3_10370: n_11751 <=  n_11752  AND n_11753  AND n_11754;
delay_10371: n_11752  <= TRANSPORT a_N1095  ;
inv_10372: n_11753  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_10373: n_11754  <= TRANSPORT dbin(3)  ;
and3_10374: n_11755 <=  n_11756  AND n_11757  AND n_11758;
delay_10375: n_11756  <= TRANSPORT a_N1095  ;
delay_10376: n_11757  <= TRANSPORT a_N2580_aNOT  ;
delay_10377: n_11758  <= TRANSPORT a_SCH3ADDRREG_F3_G  ;
and1_10378: n_11760 <=  gnd;
dff_10379: DFF_a8237

    PORT MAP ( D => a_EQ1062, CLK => a_SCH3ADDRREG_F3_G_aCLK, CLRN => a_SCH3ADDRREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F3_G);
inv_10380: a_SCH3ADDRREG_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10381: a_EQ1062 <=  n_11767  XOR n_11775;
or3_10382: n_11767 <=  n_11768  OR n_11770  OR n_11772;
and1_10383: n_11768 <=  n_11769;
delay_10384: n_11769  <= TRANSPORT a_N944_aNOT  ;
and1_10385: n_11770 <=  n_11771;
delay_10386: n_11771  <= TRANSPORT a_LC3_C26  ;
and2_10387: n_11772 <=  n_11773  AND n_11774;
delay_10388: n_11773  <= TRANSPORT a_N2528  ;
delay_10389: n_11774  <= TRANSPORT a_SCH3BAROUT_F3_G  ;
and1_10390: n_11775 <=  gnd;
delay_10391: n_11776  <= TRANSPORT clk  ;
filter_10392: FILTER_a8237

    PORT MAP (IN1 => n_11776, Y => a_SCH3ADDRREG_F3_G_aCLK);
delay_10393: a_N2544  <= TRANSPORT a_EQ601  ;
xor2_10394: a_EQ601 <=  n_11780  XOR n_11802;
or5_10395: n_11780 <=  n_11781  OR n_11785  OR n_11789  OR n_11792  OR n_11797;
and3_10396: n_11781 <=  n_11782  AND n_11783  AND n_11784;
delay_10397: n_11782  <= TRANSPORT a_N2529  ;
delay_10398: n_11783  <= TRANSPORT a_LC7_C14  ;
delay_10399: n_11784  <= TRANSPORT a_LC1_C16  ;
and3_10400: n_11785 <=  n_11786  AND n_11787  AND n_11788;
inv_10401: n_11786  <= TRANSPORT NOT a_N2529  ;
inv_10402: n_11787  <= TRANSPORT NOT a_LC7_C14  ;
delay_10403: n_11788  <= TRANSPORT a_LC1_C16  ;
and2_10404: n_11789 <=  n_11790  AND n_11791;
inv_10405: n_11790  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_10406: n_11791  <= TRANSPORT a_LC1_C16  ;
and4_10407: n_11792 <=  n_11793  AND n_11794  AND n_11795  AND n_11796;
inv_10408: n_11793  <= TRANSPORT NOT a_N2529  ;
delay_10409: n_11794  <= TRANSPORT a_N2530_aNOT  ;
delay_10410: n_11795  <= TRANSPORT a_LC7_C14  ;
inv_10411: n_11796  <= TRANSPORT NOT a_LC1_C16  ;
and4_10412: n_11797 <=  n_11798  AND n_11799  AND n_11800  AND n_11801;
delay_10413: n_11798  <= TRANSPORT a_N2529  ;
delay_10414: n_11799  <= TRANSPORT a_N2530_aNOT  ;
inv_10415: n_11800  <= TRANSPORT NOT a_LC7_C14  ;
inv_10416: n_11801  <= TRANSPORT NOT a_LC1_C16  ;
and1_10417: n_11802 <=  gnd;
delay_10418: a_LC2_C23  <= TRANSPORT a_EQ691  ;
xor2_10419: a_EQ691 <=  n_11805  XOR n_11813;
or2_10420: n_11805 <=  n_11806  OR n_11809;
and2_10421: n_11806 <=  n_11807  AND n_11808;
inv_10422: n_11807  <= TRANSPORT NOT a_N2584_aNOT  ;
delay_10423: n_11808  <= TRANSPORT dbin(4)  ;
and2_10424: n_11809 <=  n_11810  AND n_11811;
delay_10425: n_11810  <= TRANSPORT a_N2584_aNOT  ;
delay_10426: n_11811  <= TRANSPORT a_SCH1ADDRREG_F4_G  ;
and1_10427: n_11813 <=  gnd;
delay_10428: a_LC3_C23  <= TRANSPORT a_EQ692  ;
xor2_10429: a_EQ692 <=  n_11816  XOR n_11823;
or2_10430: n_11816 <=  n_11817  OR n_11820;
and2_10431: n_11817 <=  n_11818  AND n_11819;
inv_10432: n_11818  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_10433: n_11819  <= TRANSPORT a_N2544  ;
and2_10434: n_11820 <=  n_11821  AND n_11822;
delay_10435: n_11821  <= TRANSPORT a_N2559_aNOT  ;
delay_10436: n_11822  <= TRANSPORT a_LC2_C23  ;
and1_10437: n_11823 <=  gnd;
dff_10438: DFF_a8237

    PORT MAP ( D => a_EQ935, CLK => a_SCH1ADDRREG_F4_G_aCLK, CLRN => a_SCH1ADDRREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F4_G);
inv_10439: a_SCH1ADDRREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10440: a_EQ935 <=  n_11830  XOR n_11837;
or2_10441: n_11830 <=  n_11831  OR n_11834;
and2_10442: n_11831 <=  n_11832  AND n_11833;
inv_10443: n_11832  <= TRANSPORT NOT a_N2526  ;
delay_10444: n_11833  <= TRANSPORT a_LC3_C23  ;
and2_10445: n_11834 <=  n_11835  AND n_11836;
delay_10446: n_11835  <= TRANSPORT a_N2526  ;
delay_10447: n_11836  <= TRANSPORT a_SCH1BAROUT_F4_G  ;
and1_10448: n_11837 <=  gnd;
delay_10449: n_11838  <= TRANSPORT clk  ;
filter_10450: FILTER_a8237

    PORT MAP (IN1 => n_11838, Y => a_SCH1ADDRREG_F4_G_aCLK);
delay_10451: a_LC6_C5  <= TRANSPORT a_EQ287  ;
xor2_10452: a_EQ287 <=  n_11842  XOR n_11863;
or4_10453: n_11842 <=  n_11843  OR n_11848  OR n_11853  OR n_11858;
and4_10454: n_11843 <=  n_11844  AND n_11845  AND n_11846  AND n_11847;
inv_10455: n_11844  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10456: n_11845  <= TRANSPORT NOT a_N2529  ;
delay_10457: n_11846  <= TRANSPORT a_LC7_C14  ;
inv_10458: n_11847  <= TRANSPORT NOT a_LC1_C16  ;
and4_10459: n_11848 <=  n_11849  AND n_11850  AND n_11851  AND n_11852;
inv_10460: n_11849  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10461: n_11850  <= TRANSPORT a_N2529  ;
delay_10462: n_11851  <= TRANSPORT a_LC7_C14  ;
delay_10463: n_11852  <= TRANSPORT a_LC1_C16  ;
and4_10464: n_11853 <=  n_11854  AND n_11855  AND n_11856  AND n_11857;
inv_10465: n_11854  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10466: n_11855  <= TRANSPORT a_N2529  ;
inv_10467: n_11856  <= TRANSPORT NOT a_LC7_C14  ;
inv_10468: n_11857  <= TRANSPORT NOT a_LC1_C16  ;
and4_10469: n_11858 <=  n_11859  AND n_11860  AND n_11861  AND n_11862;
inv_10470: n_11859  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10471: n_11860  <= TRANSPORT NOT a_N2529  ;
inv_10472: n_11861  <= TRANSPORT NOT a_LC7_C14  ;
delay_10473: n_11862  <= TRANSPORT a_LC1_C16  ;
and1_10474: n_11863 <=  gnd;
delay_10475: a_LC3_C5  <= TRANSPORT a_EQ718  ;
xor2_10476: a_EQ718 <=  n_11866  XOR n_11876;
or2_10477: n_11866 <=  n_11867  OR n_11871;
and3_10478: n_11867 <=  n_11868  AND n_11869  AND n_11870;
delay_10479: n_11868  <= TRANSPORT a_N2560_aNOT  ;
inv_10480: n_11869  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_10481: n_11870  <= TRANSPORT dbin(4)  ;
and3_10482: n_11871 <=  n_11872  AND n_11873  AND n_11874;
delay_10483: n_11872  <= TRANSPORT a_N2560_aNOT  ;
delay_10484: n_11873  <= TRANSPORT a_N2582_aNOT  ;
delay_10485: n_11874  <= TRANSPORT a_SCH2ADDRREG_F4_G  ;
and1_10486: n_11876 <=  gnd;
dff_10487: DFF_a8237

    PORT MAP ( D => a_EQ999, CLK => a_SCH2ADDRREG_F4_G_aCLK, CLRN => a_SCH2ADDRREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F4_G);
inv_10488: a_SCH2ADDRREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10489: a_EQ999 <=  n_11883  XOR n_11893;
or3_10490: n_11883 <=  n_11884  OR n_11887  OR n_11890;
and2_10491: n_11884 <=  n_11885  AND n_11886;
inv_10492: n_11885  <= TRANSPORT NOT a_N2527  ;
delay_10493: n_11886  <= TRANSPORT a_LC6_C5  ;
and2_10494: n_11887 <=  n_11888  AND n_11889;
inv_10495: n_11888  <= TRANSPORT NOT a_N2527  ;
delay_10496: n_11889  <= TRANSPORT a_LC3_C5  ;
and2_10497: n_11890 <=  n_11891  AND n_11892;
delay_10498: n_11891  <= TRANSPORT a_N2527  ;
delay_10499: n_11892  <= TRANSPORT a_SCH2BAROUT_F4_G  ;
and1_10500: n_11893 <=  gnd;
delay_10501: n_11894  <= TRANSPORT clk  ;
filter_10502: FILTER_a8237

    PORT MAP (IN1 => n_11894, Y => a_SCH2ADDRREG_F4_G_aCLK);
delay_10503: a_N938_aNOT  <= TRANSPORT a_EQ328  ;
xor2_10504: a_EQ328 <=  n_11898  XOR n_11919;
or4_10505: n_11898 <=  n_11899  OR n_11904  OR n_11909  OR n_11914;
and4_10506: n_11899 <=  n_11900  AND n_11901  AND n_11902  AND n_11903;
delay_10507: n_11900  <= TRANSPORT a_N1094  ;
inv_10508: n_11901  <= TRANSPORT NOT a_N2529  ;
delay_10509: n_11902  <= TRANSPORT a_LC7_C14  ;
inv_10510: n_11903  <= TRANSPORT NOT a_LC1_C16  ;
and4_10511: n_11904 <=  n_11905  AND n_11906  AND n_11907  AND n_11908;
delay_10512: n_11905  <= TRANSPORT a_N1094  ;
delay_10513: n_11906  <= TRANSPORT a_N2529  ;
delay_10514: n_11907  <= TRANSPORT a_LC7_C14  ;
delay_10515: n_11908  <= TRANSPORT a_LC1_C16  ;
and4_10516: n_11909 <=  n_11910  AND n_11911  AND n_11912  AND n_11913;
delay_10517: n_11910  <= TRANSPORT a_N1094  ;
delay_10518: n_11911  <= TRANSPORT a_N2529  ;
inv_10519: n_11912  <= TRANSPORT NOT a_LC7_C14  ;
inv_10520: n_11913  <= TRANSPORT NOT a_LC1_C16  ;
and4_10521: n_11914 <=  n_11915  AND n_11916  AND n_11917  AND n_11918;
delay_10522: n_11915  <= TRANSPORT a_N1094  ;
inv_10523: n_11916  <= TRANSPORT NOT a_N2529  ;
inv_10524: n_11917  <= TRANSPORT NOT a_LC7_C14  ;
delay_10525: n_11918  <= TRANSPORT a_LC1_C16  ;
and1_10526: n_11919 <=  gnd;
delay_10527: a_LC4_C1  <= TRANSPORT a_EQ744  ;
xor2_10528: a_EQ744 <=  n_11922  XOR n_11932;
or2_10529: n_11922 <=  n_11923  OR n_11927;
and3_10530: n_11923 <=  n_11924  AND n_11925  AND n_11926;
delay_10531: n_11924  <= TRANSPORT a_N1095  ;
inv_10532: n_11925  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_10533: n_11926  <= TRANSPORT dbin(4)  ;
and3_10534: n_11927 <=  n_11928  AND n_11929  AND n_11930;
delay_10535: n_11928  <= TRANSPORT a_N1095  ;
delay_10536: n_11929  <= TRANSPORT a_N2580_aNOT  ;
delay_10537: n_11930  <= TRANSPORT a_SCH3ADDRREG_F4_G  ;
and1_10538: n_11932 <=  gnd;
dff_10539: DFF_a8237

    PORT MAP ( D => a_EQ1063, CLK => a_SCH3ADDRREG_F4_G_aCLK, CLRN => a_SCH3ADDRREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F4_G);
inv_10540: a_SCH3ADDRREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10541: a_EQ1063 <=  n_11939  XOR n_11947;
or3_10542: n_11939 <=  n_11940  OR n_11942  OR n_11944;
and1_10543: n_11940 <=  n_11941;
delay_10544: n_11941  <= TRANSPORT a_N938_aNOT  ;
and1_10545: n_11942 <=  n_11943;
delay_10546: n_11943  <= TRANSPORT a_LC4_C1  ;
and2_10547: n_11944 <=  n_11945  AND n_11946;
delay_10548: n_11945  <= TRANSPORT a_N2528  ;
delay_10549: n_11946  <= TRANSPORT a_SCH3BAROUT_F4_G  ;
and1_10550: n_11947 <=  gnd;
delay_10551: n_11948  <= TRANSPORT clk  ;
filter_10552: FILTER_a8237

    PORT MAP (IN1 => n_11948, Y => a_SCH3ADDRREG_F4_G_aCLK);
delay_10553: a_LC6_C11  <= TRANSPORT a_EQ666  ;
xor2_10554: a_EQ666 <=  n_11952  XOR n_11960;
or2_10555: n_11952 <=  n_11953  OR n_11956;
and2_10556: n_11953 <=  n_11954  AND n_11955;
delay_10557: n_11954  <= TRANSPORT a_N2586  ;
delay_10558: n_11955  <= TRANSPORT dbin(4)  ;
and2_10559: n_11956 <=  n_11957  AND n_11958;
inv_10560: n_11957  <= TRANSPORT NOT a_N2586  ;
delay_10561: n_11958  <= TRANSPORT a_SCH0ADDRREG_F4_G  ;
and1_10562: n_11960 <=  gnd;
delay_10563: a_LC5_C11  <= TRANSPORT a_EQ667  ;
xor2_10564: a_EQ667 <=  n_11963  XOR n_11970;
or2_10565: n_11963 <=  n_11964  OR n_11967;
and2_10566: n_11964 <=  n_11965  AND n_11966;
inv_10567: n_11965  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_10568: n_11966  <= TRANSPORT a_N2544  ;
and2_10569: n_11967 <=  n_11968  AND n_11969;
delay_10570: n_11968  <= TRANSPORT a_N2558_aNOT  ;
delay_10571: n_11969  <= TRANSPORT a_LC6_C11  ;
and1_10572: n_11970 <=  gnd;
dff_10573: DFF_a8237

    PORT MAP ( D => a_EQ871, CLK => a_SCH0ADDRREG_F4_G_aCLK, CLRN => a_SCH0ADDRREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F4_G);
inv_10574: a_SCH0ADDRREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10575: a_EQ871 <=  n_11977  XOR n_11984;
or2_10576: n_11977 <=  n_11978  OR n_11981;
and2_10577: n_11978 <=  n_11979  AND n_11980;
inv_10578: n_11979  <= TRANSPORT NOT a_N2525  ;
delay_10579: n_11980  <= TRANSPORT a_LC5_C11  ;
and2_10580: n_11981 <=  n_11982  AND n_11983;
delay_10581: n_11982  <= TRANSPORT a_N2525  ;
delay_10582: n_11983  <= TRANSPORT a_SCH0BAROUT_F4_G  ;
and1_10583: n_11984 <=  gnd;
delay_10584: n_11985  <= TRANSPORT clk  ;
filter_10585: FILTER_a8237

    PORT MAP (IN1 => n_11985, Y => a_SCH0ADDRREG_F4_G_aCLK);
delay_10586: a_N2545  <= TRANSPORT a_EQ602  ;
xor2_10587: a_EQ602 <=  n_11989  XOR n_12001;
or3_10588: n_11989 <=  n_11990  OR n_11994  OR n_11998;
and3_10589: n_11990 <=  n_11991  AND n_11992  AND n_11993;
inv_10590: n_11991  <= TRANSPORT NOT a_N2529  ;
delay_10591: n_11992  <= TRANSPORT a_N2530_aNOT  ;
delay_10592: n_11993  <= TRANSPORT a_LC1_F26  ;
and3_10593: n_11994 <=  n_11995  AND n_11996  AND n_11997;
delay_10594: n_11995  <= TRANSPORT a_N2529  ;
delay_10595: n_11996  <= TRANSPORT a_N2530_aNOT  ;
inv_10596: n_11997  <= TRANSPORT NOT a_LC1_F26  ;
and2_10597: n_11998 <=  n_11999  AND n_12000;
inv_10598: n_11999  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_10599: n_12000  <= TRANSPORT a_LC3_F6  ;
and1_10600: n_12001 <=  gnd;
delay_10601: a_LC2_F23  <= TRANSPORT a_EQ689  ;
xor2_10602: a_EQ689 <=  n_12004  XOR n_12016;
or3_10603: n_12004 <=  n_12005  OR n_12009  OR n_12012;
and2_10604: n_12005 <=  n_12006  AND n_12007;
delay_10605: n_12006  <= TRANSPORT a_N2352  ;
delay_10606: n_12007  <= TRANSPORT a_SCH1ADDRREG_F5_G  ;
and2_10607: n_12009 <=  n_12010  AND n_12011;
delay_10608: n_12010  <= TRANSPORT a_LC6_D6  ;
delay_10609: n_12011  <= TRANSPORT a_SCH1ADDRREG_F5_G  ;
and3_10610: n_12012 <=  n_12013  AND n_12014  AND n_12015;
inv_10611: n_12013  <= TRANSPORT NOT a_LC6_D6  ;
inv_10612: n_12014  <= TRANSPORT NOT a_N2352  ;
delay_10613: n_12015  <= TRANSPORT dbin(5)  ;
and1_10614: n_12016 <=  gnd;
delay_10615: a_LC4_F23  <= TRANSPORT a_EQ690  ;
xor2_10616: a_EQ690 <=  n_12019  XOR n_12026;
or2_10617: n_12019 <=  n_12020  OR n_12023;
and2_10618: n_12020 <=  n_12021  AND n_12022;
inv_10619: n_12021  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_10620: n_12022  <= TRANSPORT a_N2545  ;
and2_10621: n_12023 <=  n_12024  AND n_12025;
delay_10622: n_12024  <= TRANSPORT a_N2559_aNOT  ;
delay_10623: n_12025  <= TRANSPORT a_LC2_F23  ;
and1_10624: n_12026 <=  gnd;
dff_10625: DFF_a8237

    PORT MAP ( D => a_EQ936, CLK => a_SCH1ADDRREG_F5_G_aCLK, CLRN => a_SCH1ADDRREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F5_G);
inv_10626: a_SCH1ADDRREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10627: a_EQ936 <=  n_12033  XOR n_12044;
or3_10628: n_12033 <=  n_12034  OR n_12037  OR n_12040;
and2_10629: n_12034 <=  n_12035  AND n_12036;
inv_10630: n_12035  <= TRANSPORT NOT a_SCH1MODEREG_F2_G  ;
delay_10631: n_12036  <= TRANSPORT a_LC4_F23  ;
and2_10632: n_12037 <=  n_12038  AND n_12039;
inv_10633: n_12038  <= TRANSPORT NOT a_N57_aNOT  ;
delay_10634: n_12039  <= TRANSPORT a_LC4_F23  ;
and3_10635: n_12040 <=  n_12041  AND n_12042  AND n_12043;
delay_10636: n_12041  <= TRANSPORT a_N57_aNOT  ;
delay_10637: n_12042  <= TRANSPORT a_SCH1BAROUT_F5_G  ;
delay_10638: n_12043  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and1_10639: n_12044 <=  gnd;
delay_10640: n_12045  <= TRANSPORT clk  ;
filter_10641: FILTER_a8237

    PORT MAP (IN1 => n_12045, Y => a_SCH1ADDRREG_F5_G_aCLK);
delay_10642: a_LC3_F20  <= TRANSPORT a_EQ716  ;
xor2_10643: a_EQ716 <=  n_12049  XOR n_12057;
or2_10644: n_12049 <=  n_12050  OR n_12053;
and2_10645: n_12050 <=  n_12051  AND n_12052;
inv_10646: n_12051  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_10647: n_12052  <= TRANSPORT dbin(5)  ;
and2_10648: n_12053 <=  n_12054  AND n_12055;
delay_10649: n_12054  <= TRANSPORT a_N2582_aNOT  ;
delay_10650: n_12055  <= TRANSPORT a_SCH2ADDRREG_F5_G  ;
and1_10651: n_12057 <=  gnd;
delay_10652: a_LC1_F20  <= TRANSPORT a_EQ717  ;
xor2_10653: a_EQ717 <=  n_12060  XOR n_12072;
or3_10654: n_12060 <=  n_12061  OR n_12065  OR n_12069;
and3_10655: n_12061 <=  n_12062  AND n_12063  AND n_12064;
inv_10656: n_12062  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10657: n_12063  <= TRANSPORT NOT a_N2529  ;
delay_10658: n_12064  <= TRANSPORT a_LC1_F26  ;
and3_10659: n_12065 <=  n_12066  AND n_12067  AND n_12068;
inv_10660: n_12066  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10661: n_12067  <= TRANSPORT a_N2529  ;
inv_10662: n_12068  <= TRANSPORT NOT a_LC1_F26  ;
and2_10663: n_12069 <=  n_12070  AND n_12071;
delay_10664: n_12070  <= TRANSPORT a_N2560_aNOT  ;
delay_10665: n_12071  <= TRANSPORT a_LC3_F20  ;
and1_10666: n_12072 <=  gnd;
dff_10667: DFF_a8237

    PORT MAP ( D => a_EQ1000, CLK => a_SCH2ADDRREG_F5_G_aCLK, CLRN => a_SCH2ADDRREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F5_G);
inv_10668: a_SCH2ADDRREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10669: a_EQ1000 <=  n_12079  XOR n_12086;
or2_10670: n_12079 <=  n_12080  OR n_12083;
and2_10671: n_12080 <=  n_12081  AND n_12082;
inv_10672: n_12081  <= TRANSPORT NOT a_N2527  ;
delay_10673: n_12082  <= TRANSPORT a_LC1_F20  ;
and2_10674: n_12083 <=  n_12084  AND n_12085;
delay_10675: n_12084  <= TRANSPORT a_N2527  ;
delay_10676: n_12085  <= TRANSPORT a_SCH2BAROUT_F5_G  ;
and1_10677: n_12086 <=  gnd;
delay_10678: n_12087  <= TRANSPORT clk  ;
filter_10679: FILTER_a8237

    PORT MAP (IN1 => n_12087, Y => a_SCH2ADDRREG_F5_G_aCLK);
delay_10680: a_LC1_F21  <= TRANSPORT a_EQ742  ;
xor2_10681: a_EQ742 <=  n_12091  XOR n_12101;
or2_10682: n_12091 <=  n_12092  OR n_12096;
and3_10683: n_12092 <=  n_12093  AND n_12094  AND n_12095;
delay_10684: n_12093  <= TRANSPORT a_N1095  ;
inv_10685: n_12094  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_10686: n_12095  <= TRANSPORT dbin(5)  ;
and3_10687: n_12096 <=  n_12097  AND n_12098  AND n_12099;
delay_10688: n_12097  <= TRANSPORT a_N1095  ;
delay_10689: n_12098  <= TRANSPORT a_N2580_aNOT  ;
delay_10690: n_12099  <= TRANSPORT a_SCH3ADDRREG_F5_G  ;
and1_10691: n_12101 <=  gnd;
delay_10692: a_LC3_F21  <= TRANSPORT a_EQ743  ;
xor2_10693: a_EQ743 <=  n_12104  XOR n_12110;
or2_10694: n_12104 <=  n_12105  OR n_12107;
and1_10695: n_12105 <=  n_12106;
delay_10696: n_12106  <= TRANSPORT a_LC1_F21  ;
and2_10697: n_12107 <=  n_12108  AND n_12109;
delay_10698: n_12108  <= TRANSPORT a_N2528  ;
delay_10699: n_12109  <= TRANSPORT a_SCH3BAROUT_F5_G  ;
and1_10700: n_12110 <=  gnd;
dff_10701: DFF_a8237

    PORT MAP ( D => a_EQ1064, CLK => a_SCH3ADDRREG_F5_G_aCLK, CLRN => a_SCH3ADDRREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F5_G);
inv_10702: a_SCH3ADDRREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10703: a_EQ1064 <=  n_12117  XOR n_12128;
or3_10704: n_12117 <=  n_12118  OR n_12120  OR n_12124;
and1_10705: n_12118 <=  n_12119;
delay_10706: n_12119  <= TRANSPORT a_LC3_F21  ;
and3_10707: n_12120 <=  n_12121  AND n_12122  AND n_12123;
delay_10708: n_12121  <= TRANSPORT a_N1094  ;
inv_10709: n_12122  <= TRANSPORT NOT a_N2529  ;
delay_10710: n_12123  <= TRANSPORT a_LC1_F26  ;
and3_10711: n_12124 <=  n_12125  AND n_12126  AND n_12127;
delay_10712: n_12125  <= TRANSPORT a_N1094  ;
delay_10713: n_12126  <= TRANSPORT a_N2529  ;
inv_10714: n_12127  <= TRANSPORT NOT a_LC1_F26  ;
and1_10715: n_12128 <=  gnd;
delay_10716: n_12129  <= TRANSPORT clk  ;
filter_10717: FILTER_a8237

    PORT MAP (IN1 => n_12129, Y => a_SCH3ADDRREG_F5_G_aCLK);
delay_10718: a_LC3_F3  <= TRANSPORT a_EQ664  ;
xor2_10719: a_EQ664 <=  n_12133  XOR n_12145;
or3_10720: n_12133 <=  n_12134  OR n_12138  OR n_12141;
and2_10721: n_12134 <=  n_12135  AND n_12136;
inv_10722: n_12135  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_10723: n_12136  <= TRANSPORT a_SCH0ADDRREG_F5_G  ;
and2_10724: n_12138 <=  n_12139  AND n_12140;
delay_10725: n_12139  <= TRANSPORT a_LC6_D6  ;
delay_10726: n_12140  <= TRANSPORT a_SCH0ADDRREG_F5_G  ;
and3_10727: n_12141 <=  n_12142  AND n_12143  AND n_12144;
inv_10728: n_12142  <= TRANSPORT NOT a_LC6_D6  ;
delay_10729: n_12143  <= TRANSPORT a_N2354_aNOT  ;
delay_10730: n_12144  <= TRANSPORT dbin(5)  ;
and1_10731: n_12145 <=  gnd;
delay_10732: a_LC4_F3  <= TRANSPORT a_EQ665  ;
xor2_10733: a_EQ665 <=  n_12148  XOR n_12155;
or2_10734: n_12148 <=  n_12149  OR n_12152;
and2_10735: n_12149 <=  n_12150  AND n_12151;
inv_10736: n_12150  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_10737: n_12151  <= TRANSPORT a_N2545  ;
and2_10738: n_12152 <=  n_12153  AND n_12154;
delay_10739: n_12153  <= TRANSPORT a_N2558_aNOT  ;
delay_10740: n_12154  <= TRANSPORT a_LC3_F3  ;
and1_10741: n_12155 <=  gnd;
dff_10742: DFF_a8237

    PORT MAP ( D => a_EQ872, CLK => a_SCH0ADDRREG_F5_G_aCLK, CLRN => a_SCH0ADDRREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F5_G);
inv_10743: a_SCH0ADDRREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10744: a_EQ872 <=  n_12162  XOR n_12173;
or3_10745: n_12162 <=  n_12163  OR n_12166  OR n_12169;
and2_10746: n_12163 <=  n_12164  AND n_12165;
inv_10747: n_12164  <= TRANSPORT NOT a_SCH0MODEREG_F2_G  ;
delay_10748: n_12165  <= TRANSPORT a_LC4_F3  ;
and2_10749: n_12166 <=  n_12167  AND n_12168;
inv_10750: n_12167  <= TRANSPORT NOT a_N57_aNOT  ;
delay_10751: n_12168  <= TRANSPORT a_LC4_F3  ;
and3_10752: n_12169 <=  n_12170  AND n_12171  AND n_12172;
delay_10753: n_12170  <= TRANSPORT a_N57_aNOT  ;
delay_10754: n_12171  <= TRANSPORT a_SCH0BAROUT_F5_G  ;
delay_10755: n_12172  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and1_10756: n_12173 <=  gnd;
delay_10757: n_12174  <= TRANSPORT clk  ;
filter_10758: FILTER_a8237

    PORT MAP (IN1 => n_12174, Y => a_SCH0ADDRREG_F5_G_aCLK);
delay_10759: a_LC3_F14  <= TRANSPORT a_EQ288  ;
xor2_10760: a_EQ288 <=  n_12178  XOR n_12199;
or4_10761: n_12178 <=  n_12179  OR n_12184  OR n_12189  OR n_12194;
and4_10762: n_12179 <=  n_12180  AND n_12181  AND n_12182  AND n_12183;
inv_10763: n_12180  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10764: n_12181  <= TRANSPORT NOT a_N2529  ;
delay_10765: n_12182  <= TRANSPORT a_LC6_F20  ;
inv_10766: n_12183  <= TRANSPORT NOT a_LC4_F10  ;
and4_10767: n_12184 <=  n_12185  AND n_12186  AND n_12187  AND n_12188;
inv_10768: n_12185  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10769: n_12186  <= TRANSPORT a_N2529  ;
delay_10770: n_12187  <= TRANSPORT a_LC6_F20  ;
delay_10771: n_12188  <= TRANSPORT a_LC4_F10  ;
and4_10772: n_12189 <=  n_12190  AND n_12191  AND n_12192  AND n_12193;
inv_10773: n_12190  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_10774: n_12191  <= TRANSPORT a_N2529  ;
inv_10775: n_12192  <= TRANSPORT NOT a_LC6_F20  ;
inv_10776: n_12193  <= TRANSPORT NOT a_LC4_F10  ;
and4_10777: n_12194 <=  n_12195  AND n_12196  AND n_12197  AND n_12198;
inv_10778: n_12195  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_10779: n_12196  <= TRANSPORT NOT a_N2529  ;
inv_10780: n_12197  <= TRANSPORT NOT a_LC6_F20  ;
delay_10781: n_12198  <= TRANSPORT a_LC4_F10  ;
and1_10782: n_12199 <=  gnd;
delay_10783: a_LC4_F14  <= TRANSPORT a_EQ715  ;
xor2_10784: a_EQ715 <=  n_12202  XOR n_12212;
or2_10785: n_12202 <=  n_12203  OR n_12207;
and3_10786: n_12203 <=  n_12204  AND n_12205  AND n_12206;
delay_10787: n_12204  <= TRANSPORT a_N2560_aNOT  ;
inv_10788: n_12205  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_10789: n_12206  <= TRANSPORT dbin(6)  ;
and3_10790: n_12207 <=  n_12208  AND n_12209  AND n_12210;
delay_10791: n_12208  <= TRANSPORT a_N2560_aNOT  ;
delay_10792: n_12209  <= TRANSPORT a_N2582_aNOT  ;
delay_10793: n_12210  <= TRANSPORT a_SCH2ADDRREG_F6_G  ;
and1_10794: n_12212 <=  gnd;
dff_10795: DFF_a8237

    PORT MAP ( D => a_EQ1001, CLK => a_SCH2ADDRREG_F6_G_aCLK, CLRN => a_SCH2ADDRREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F6_G);
inv_10796: a_SCH2ADDRREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10797: a_EQ1001 <=  n_12219  XOR n_12229;
or3_10798: n_12219 <=  n_12220  OR n_12223  OR n_12226;
and2_10799: n_12220 <=  n_12221  AND n_12222;
inv_10800: n_12221  <= TRANSPORT NOT a_N2527  ;
delay_10801: n_12222  <= TRANSPORT a_LC3_F14  ;
and2_10802: n_12223 <=  n_12224  AND n_12225;
inv_10803: n_12224  <= TRANSPORT NOT a_N2527  ;
delay_10804: n_12225  <= TRANSPORT a_LC4_F14  ;
and2_10805: n_12226 <=  n_12227  AND n_12228;
delay_10806: n_12227  <= TRANSPORT a_N2527  ;
delay_10807: n_12228  <= TRANSPORT a_SCH2BAROUT_F6_G  ;
and1_10808: n_12229 <=  gnd;
delay_10809: n_12230  <= TRANSPORT clk  ;
filter_10810: FILTER_a8237

    PORT MAP (IN1 => n_12230, Y => a_SCH2ADDRREG_F6_G_aCLK);
delay_10811: a_N2546  <= TRANSPORT a_EQ603  ;
xor2_10812: a_EQ603 <=  n_12234  XOR n_12256;
or5_10813: n_12234 <=  n_12235  OR n_12239  OR n_12243  OR n_12246  OR n_12251;
and3_10814: n_12235 <=  n_12236  AND n_12237  AND n_12238;
delay_10815: n_12236  <= TRANSPORT a_N2529  ;
delay_10816: n_12237  <= TRANSPORT a_LC6_F20  ;
delay_10817: n_12238  <= TRANSPORT a_LC4_F10  ;
and3_10818: n_12239 <=  n_12240  AND n_12241  AND n_12242;
inv_10819: n_12240  <= TRANSPORT NOT a_N2529  ;
inv_10820: n_12241  <= TRANSPORT NOT a_LC6_F20  ;
delay_10821: n_12242  <= TRANSPORT a_LC4_F10  ;
and2_10822: n_12243 <=  n_12244  AND n_12245;
inv_10823: n_12244  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_10824: n_12245  <= TRANSPORT a_LC4_F10  ;
and4_10825: n_12246 <=  n_12247  AND n_12248  AND n_12249  AND n_12250;
inv_10826: n_12247  <= TRANSPORT NOT a_N2529  ;
delay_10827: n_12248  <= TRANSPORT a_N2530_aNOT  ;
delay_10828: n_12249  <= TRANSPORT a_LC6_F20  ;
inv_10829: n_12250  <= TRANSPORT NOT a_LC4_F10  ;
and4_10830: n_12251 <=  n_12252  AND n_12253  AND n_12254  AND n_12255;
delay_10831: n_12252  <= TRANSPORT a_N2529  ;
delay_10832: n_12253  <= TRANSPORT a_N2530_aNOT  ;
inv_10833: n_12254  <= TRANSPORT NOT a_LC6_F20  ;
inv_10834: n_12255  <= TRANSPORT NOT a_LC4_F10  ;
and1_10835: n_12256 <=  gnd;
delay_10836: a_LC5_F3  <= TRANSPORT a_EQ662  ;
xor2_10837: a_EQ662 <=  n_12259  XOR n_12271;
or3_10838: n_12259 <=  n_12260  OR n_12264  OR n_12267;
and2_10839: n_12260 <=  n_12261  AND n_12262;
inv_10840: n_12261  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_10841: n_12262  <= TRANSPORT a_SCH0ADDRREG_F6_G  ;
and2_10842: n_12264 <=  n_12265  AND n_12266;
delay_10843: n_12265  <= TRANSPORT a_LC6_D6  ;
delay_10844: n_12266  <= TRANSPORT a_SCH0ADDRREG_F6_G  ;
and3_10845: n_12267 <=  n_12268  AND n_12269  AND n_12270;
inv_10846: n_12268  <= TRANSPORT NOT a_LC6_D6  ;
delay_10847: n_12269  <= TRANSPORT a_N2354_aNOT  ;
delay_10848: n_12270  <= TRANSPORT dbin(6)  ;
and1_10849: n_12271 <=  gnd;
delay_10850: a_LC2_F3  <= TRANSPORT a_EQ663  ;
xor2_10851: a_EQ663 <=  n_12274  XOR n_12281;
or2_10852: n_12274 <=  n_12275  OR n_12278;
and2_10853: n_12275 <=  n_12276  AND n_12277;
inv_10854: n_12276  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_10855: n_12277  <= TRANSPORT a_N2546  ;
and2_10856: n_12278 <=  n_12279  AND n_12280;
delay_10857: n_12279  <= TRANSPORT a_N2558_aNOT  ;
delay_10858: n_12280  <= TRANSPORT a_LC5_F3  ;
and1_10859: n_12281 <=  gnd;
dff_10860: DFF_a8237

    PORT MAP ( D => a_EQ873, CLK => a_SCH0ADDRREG_F6_G_aCLK, CLRN => a_SCH0ADDRREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F6_G);
inv_10861: a_SCH0ADDRREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10862: a_EQ873 <=  n_12288  XOR n_12299;
or3_10863: n_12288 <=  n_12289  OR n_12292  OR n_12295;
and2_10864: n_12289 <=  n_12290  AND n_12291;
inv_10865: n_12290  <= TRANSPORT NOT a_SCH0MODEREG_F2_G  ;
delay_10866: n_12291  <= TRANSPORT a_LC2_F3  ;
and2_10867: n_12292 <=  n_12293  AND n_12294;
inv_10868: n_12293  <= TRANSPORT NOT a_N57_aNOT  ;
delay_10869: n_12294  <= TRANSPORT a_LC2_F3  ;
and3_10870: n_12295 <=  n_12296  AND n_12297  AND n_12298;
delay_10871: n_12296  <= TRANSPORT a_N57_aNOT  ;
delay_10872: n_12297  <= TRANSPORT a_SCH0BAROUT_F6_G  ;
delay_10873: n_12298  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and1_10874: n_12299 <=  gnd;
delay_10875: n_12300  <= TRANSPORT clk  ;
filter_10876: FILTER_a8237

    PORT MAP (IN1 => n_12300, Y => a_SCH0ADDRREG_F6_G_aCLK);
delay_10877: a_LC5_F23  <= TRANSPORT a_EQ687  ;
xor2_10878: a_EQ687 <=  n_12304  XOR n_12316;
or3_10879: n_12304 <=  n_12305  OR n_12309  OR n_12312;
and2_10880: n_12305 <=  n_12306  AND n_12307;
delay_10881: n_12306  <= TRANSPORT a_N2352  ;
delay_10882: n_12307  <= TRANSPORT a_SCH1ADDRREG_F6_G  ;
and2_10883: n_12309 <=  n_12310  AND n_12311;
delay_10884: n_12310  <= TRANSPORT a_LC6_D6  ;
delay_10885: n_12311  <= TRANSPORT a_SCH1ADDRREG_F6_G  ;
and3_10886: n_12312 <=  n_12313  AND n_12314  AND n_12315;
inv_10887: n_12313  <= TRANSPORT NOT a_LC6_D6  ;
inv_10888: n_12314  <= TRANSPORT NOT a_N2352  ;
delay_10889: n_12315  <= TRANSPORT dbin(6)  ;
and1_10890: n_12316 <=  gnd;
delay_10891: a_LC1_F23  <= TRANSPORT a_EQ688  ;
xor2_10892: a_EQ688 <=  n_12319  XOR n_12326;
or2_10893: n_12319 <=  n_12320  OR n_12323;
and2_10894: n_12320 <=  n_12321  AND n_12322;
inv_10895: n_12321  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_10896: n_12322  <= TRANSPORT a_N2546  ;
and2_10897: n_12323 <=  n_12324  AND n_12325;
delay_10898: n_12324  <= TRANSPORT a_N2559_aNOT  ;
delay_10899: n_12325  <= TRANSPORT a_LC5_F23  ;
and1_10900: n_12326 <=  gnd;
dff_10901: DFF_a8237

    PORT MAP ( D => a_EQ937, CLK => a_SCH1ADDRREG_F6_G_aCLK, CLRN => a_SCH1ADDRREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F6_G);
inv_10902: a_SCH1ADDRREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10903: a_EQ937 <=  n_12333  XOR n_12344;
or3_10904: n_12333 <=  n_12334  OR n_12337  OR n_12340;
and2_10905: n_12334 <=  n_12335  AND n_12336;
inv_10906: n_12335  <= TRANSPORT NOT a_SCH1MODEREG_F2_G  ;
delay_10907: n_12336  <= TRANSPORT a_LC1_F23  ;
and2_10908: n_12337 <=  n_12338  AND n_12339;
inv_10909: n_12338  <= TRANSPORT NOT a_N57_aNOT  ;
delay_10910: n_12339  <= TRANSPORT a_LC1_F23  ;
and3_10911: n_12340 <=  n_12341  AND n_12342  AND n_12343;
delay_10912: n_12341  <= TRANSPORT a_N57_aNOT  ;
delay_10913: n_12342  <= TRANSPORT a_SCH1BAROUT_F6_G  ;
delay_10914: n_12343  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and1_10915: n_12344 <=  gnd;
delay_10916: n_12345  <= TRANSPORT clk  ;
filter_10917: FILTER_a8237

    PORT MAP (IN1 => n_12345, Y => a_SCH1ADDRREG_F6_G_aCLK);
delay_10918: a_N933_aNOT  <= TRANSPORT a_EQ326  ;
xor2_10919: a_EQ326 <=  n_12349  XOR n_12370;
or4_10920: n_12349 <=  n_12350  OR n_12355  OR n_12360  OR n_12365;
and4_10921: n_12350 <=  n_12351  AND n_12352  AND n_12353  AND n_12354;
delay_10922: n_12351  <= TRANSPORT a_N1094  ;
inv_10923: n_12352  <= TRANSPORT NOT a_N2529  ;
delay_10924: n_12353  <= TRANSPORT a_LC6_F20  ;
inv_10925: n_12354  <= TRANSPORT NOT a_LC4_F10  ;
and4_10926: n_12355 <=  n_12356  AND n_12357  AND n_12358  AND n_12359;
delay_10927: n_12356  <= TRANSPORT a_N1094  ;
delay_10928: n_12357  <= TRANSPORT a_N2529  ;
delay_10929: n_12358  <= TRANSPORT a_LC6_F20  ;
delay_10930: n_12359  <= TRANSPORT a_LC4_F10  ;
and4_10931: n_12360 <=  n_12361  AND n_12362  AND n_12363  AND n_12364;
delay_10932: n_12361  <= TRANSPORT a_N1094  ;
delay_10933: n_12362  <= TRANSPORT a_N2529  ;
inv_10934: n_12363  <= TRANSPORT NOT a_LC6_F20  ;
inv_10935: n_12364  <= TRANSPORT NOT a_LC4_F10  ;
and4_10936: n_12365 <=  n_12366  AND n_12367  AND n_12368  AND n_12369;
delay_10937: n_12366  <= TRANSPORT a_N1094  ;
inv_10938: n_12367  <= TRANSPORT NOT a_N2529  ;
inv_10939: n_12368  <= TRANSPORT NOT a_LC6_F20  ;
delay_10940: n_12369  <= TRANSPORT a_LC4_F10  ;
and1_10941: n_12370 <=  gnd;
delay_10942: a_LC4_F21  <= TRANSPORT a_EQ741  ;
xor2_10943: a_EQ741 <=  n_12373  XOR n_12383;
or2_10944: n_12373 <=  n_12374  OR n_12378;
and3_10945: n_12374 <=  n_12375  AND n_12376  AND n_12377;
delay_10946: n_12375  <= TRANSPORT a_N1095  ;
inv_10947: n_12376  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_10948: n_12377  <= TRANSPORT dbin(6)  ;
and3_10949: n_12378 <=  n_12379  AND n_12380  AND n_12381;
delay_10950: n_12379  <= TRANSPORT a_N1095  ;
delay_10951: n_12380  <= TRANSPORT a_N2580_aNOT  ;
delay_10952: n_12381  <= TRANSPORT a_SCH3ADDRREG_F6_G  ;
and1_10953: n_12383 <=  gnd;
dff_10954: DFF_a8237

    PORT MAP ( D => a_EQ1065, CLK => a_SCH3ADDRREG_F6_G_aCLK, CLRN => a_SCH3ADDRREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F6_G);
inv_10955: a_SCH3ADDRREG_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10956: a_EQ1065 <=  n_12390  XOR n_12398;
or3_10957: n_12390 <=  n_12391  OR n_12393  OR n_12395;
and1_10958: n_12391 <=  n_12392;
delay_10959: n_12392  <= TRANSPORT a_N933_aNOT  ;
and1_10960: n_12393 <=  n_12394;
delay_10961: n_12394  <= TRANSPORT a_LC4_F21  ;
and2_10962: n_12395 <=  n_12396  AND n_12397;
delay_10963: n_12396  <= TRANSPORT a_N2528  ;
delay_10964: n_12397  <= TRANSPORT a_SCH3BAROUT_F6_G  ;
and1_10965: n_12398 <=  gnd;
delay_10966: n_12399  <= TRANSPORT clk  ;
filter_10967: FILTER_a8237

    PORT MAP (IN1 => n_12399, Y => a_SCH3ADDRREG_F6_G_aCLK);
delay_10968: a_LC6_D25  <= TRANSPORT a_EQ739  ;
xor2_10969: a_EQ739 <=  n_12403  XOR n_12413;
or2_10970: n_12403 <=  n_12404  OR n_12408;
and3_10971: n_12404 <=  n_12405  AND n_12406  AND n_12407;
delay_10972: n_12405  <= TRANSPORT a_N1095  ;
inv_10973: n_12406  <= TRANSPORT NOT a_N2580_aNOT  ;
delay_10974: n_12407  <= TRANSPORT dbin(7)  ;
and3_10975: n_12408 <=  n_12409  AND n_12410  AND n_12411;
delay_10976: n_12409  <= TRANSPORT a_N1095  ;
delay_10977: n_12410  <= TRANSPORT a_N2580_aNOT  ;
delay_10978: n_12411  <= TRANSPORT a_SCH3ADDRREG_F7_G  ;
and1_10979: n_12413 <=  gnd;
delay_10980: a_LC4_D25  <= TRANSPORT a_EQ740  ;
xor2_10981: a_EQ740 <=  n_12416  XOR n_12422;
or2_10982: n_12416 <=  n_12417  OR n_12419;
and1_10983: n_12417 <=  n_12418;
delay_10984: n_12418  <= TRANSPORT a_LC6_D25  ;
and2_10985: n_12419 <=  n_12420  AND n_12421;
delay_10986: n_12420  <= TRANSPORT a_N2528  ;
delay_10987: n_12421  <= TRANSPORT a_SCH3BAROUT_F7_G  ;
and1_10988: n_12422 <=  gnd;
dff_10989: DFF_a8237

    PORT MAP ( D => a_EQ1066, CLK => a_SCH3ADDRREG_F7_G_aCLK, CLRN => a_SCH3ADDRREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH3ADDRREG_F7_G);
inv_10990: a_SCH3ADDRREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_10991: a_EQ1066 <=  n_12429  XOR n_12440;
or3_10992: n_12429 <=  n_12430  OR n_12434  OR n_12438;
and3_10993: n_12430 <=  n_12431  AND n_12432  AND n_12433;
delay_10994: n_12431  <= TRANSPORT a_N1094  ;
inv_10995: n_12432  <= TRANSPORT NOT a_N2529  ;
delay_10996: n_12433  <= TRANSPORT a_LC4_F15  ;
and3_10997: n_12434 <=  n_12435  AND n_12436  AND n_12437;
delay_10998: n_12435  <= TRANSPORT a_N1094  ;
delay_10999: n_12436  <= TRANSPORT a_N2529  ;
inv_11000: n_12437  <= TRANSPORT NOT a_LC4_F15  ;
and1_11001: n_12438 <=  n_12439;
delay_11002: n_12439  <= TRANSPORT a_LC4_D25  ;
and1_11003: n_12440 <=  gnd;
delay_11004: n_12441  <= TRANSPORT clk  ;
filter_11005: FILTER_a8237

    PORT MAP (IN1 => n_12441, Y => a_SCH3ADDRREG_F7_G_aCLK);
delay_11006: a_N786_aNOT  <= TRANSPORT a_EQ299  ;
xor2_11007: a_EQ299 <=  n_12445  XOR n_12453;
or2_11008: n_12445 <=  n_12446  OR n_12449;
and2_11009: n_12446 <=  n_12447  AND n_12448;
inv_11010: n_12447  <= TRANSPORT NOT a_N2582_aNOT  ;
delay_11011: n_12448  <= TRANSPORT dbin(7)  ;
and2_11012: n_12449 <=  n_12450  AND n_12451;
delay_11013: n_12450  <= TRANSPORT a_N2582_aNOT  ;
delay_11014: n_12451  <= TRANSPORT a_SCH2ADDRREG_F7_G  ;
and1_11015: n_12453 <=  gnd;
delay_11016: a_LC4_D17  <= TRANSPORT a_EQ714  ;
xor2_11017: a_EQ714 <=  n_12456  XOR n_12468;
or3_11018: n_12456 <=  n_12457  OR n_12461  OR n_12465;
and3_11019: n_12457 <=  n_12458  AND n_12459  AND n_12460;
inv_11020: n_12458  <= TRANSPORT NOT a_N2560_aNOT  ;
inv_11021: n_12459  <= TRANSPORT NOT a_N2529  ;
delay_11022: n_12460  <= TRANSPORT a_LC4_F15  ;
and3_11023: n_12461 <=  n_12462  AND n_12463  AND n_12464;
inv_11024: n_12462  <= TRANSPORT NOT a_N2560_aNOT  ;
delay_11025: n_12463  <= TRANSPORT a_N2529  ;
inv_11026: n_12464  <= TRANSPORT NOT a_LC4_F15  ;
and2_11027: n_12465 <=  n_12466  AND n_12467;
delay_11028: n_12466  <= TRANSPORT a_N2560_aNOT  ;
delay_11029: n_12467  <= TRANSPORT a_N786_aNOT  ;
and1_11030: n_12468 <=  gnd;
dff_11031: DFF_a8237

    PORT MAP ( D => a_EQ1002, CLK => a_SCH2ADDRREG_F7_G_aCLK, CLRN => a_SCH2ADDRREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH2ADDRREG_F7_G);
inv_11032: a_SCH2ADDRREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11033: a_EQ1002 <=  n_12475  XOR n_12482;
or2_11034: n_12475 <=  n_12476  OR n_12479;
and2_11035: n_12476 <=  n_12477  AND n_12478;
inv_11036: n_12477  <= TRANSPORT NOT a_N2527  ;
delay_11037: n_12478  <= TRANSPORT a_LC4_D17  ;
and2_11038: n_12479 <=  n_12480  AND n_12481;
delay_11039: n_12480  <= TRANSPORT a_N2527  ;
delay_11040: n_12481  <= TRANSPORT a_SCH2BAROUT_F7_G  ;
and1_11041: n_12482 <=  gnd;
delay_11042: n_12483  <= TRANSPORT clk  ;
filter_11043: FILTER_a8237

    PORT MAP (IN1 => n_12483, Y => a_SCH2ADDRREG_F7_G_aCLK);
delay_11044: a_N2547  <= TRANSPORT a_EQ604  ;
xor2_11045: a_EQ604 <=  n_12487  XOR n_12509;
or5_11046: n_12487 <=  n_12488  OR n_12492  OR n_12496  OR n_12499  OR n_12504;
and3_11047: n_12488 <=  n_12489  AND n_12490  AND n_12491;
delay_11048: n_12489  <= TRANSPORT a_N2529  ;
delay_11049: n_12490  <= TRANSPORT a_LC6_F15  ;
delay_11050: n_12491  <= TRANSPORT a_LC5_D27  ;
and3_11051: n_12492 <=  n_12493  AND n_12494  AND n_12495;
inv_11052: n_12493  <= TRANSPORT NOT a_N2529  ;
inv_11053: n_12494  <= TRANSPORT NOT a_LC6_F15  ;
delay_11054: n_12495  <= TRANSPORT a_LC5_D27  ;
and2_11055: n_12496 <=  n_12497  AND n_12498;
inv_11056: n_12497  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_11057: n_12498  <= TRANSPORT a_LC5_D27  ;
and4_11058: n_12499 <=  n_12500  AND n_12501  AND n_12502  AND n_12503;
inv_11059: n_12500  <= TRANSPORT NOT a_N2529  ;
delay_11060: n_12501  <= TRANSPORT a_N2530_aNOT  ;
delay_11061: n_12502  <= TRANSPORT a_LC6_F15  ;
inv_11062: n_12503  <= TRANSPORT NOT a_LC5_D27  ;
and4_11063: n_12504 <=  n_12505  AND n_12506  AND n_12507  AND n_12508;
delay_11064: n_12505  <= TRANSPORT a_N2529  ;
delay_11065: n_12506  <= TRANSPORT a_N2530_aNOT  ;
inv_11066: n_12507  <= TRANSPORT NOT a_LC6_F15  ;
inv_11067: n_12508  <= TRANSPORT NOT a_LC5_D27  ;
and1_11068: n_12509 <=  gnd;
delay_11069: a_N183_aNOT  <= TRANSPORT a_EQ204  ;
xor2_11070: a_EQ204 <=  n_12512  XOR n_12524;
or3_11071: n_12512 <=  n_12513  OR n_12517  OR n_12521;
and3_11072: n_12513 <=  n_12514  AND n_12515  AND n_12516;
inv_11073: n_12514  <= TRANSPORT NOT a_LC6_D6  ;
delay_11074: n_12515  <= TRANSPORT a_N2354_aNOT  ;
delay_11075: n_12516  <= TRANSPORT dbin(7)  ;
and2_11076: n_12517 <=  n_12518  AND n_12519;
inv_11077: n_12518  <= TRANSPORT NOT a_N2354_aNOT  ;
delay_11078: n_12519  <= TRANSPORT a_SCH0ADDRREG_F7_G  ;
and2_11079: n_12521 <=  n_12522  AND n_12523;
delay_11080: n_12522  <= TRANSPORT a_LC6_D6  ;
delay_11081: n_12523  <= TRANSPORT a_SCH0ADDRREG_F7_G  ;
and1_11082: n_12524 <=  gnd;
delay_11083: a_LC3_D9  <= TRANSPORT a_EQ661  ;
xor2_11084: a_EQ661 <=  n_12527  XOR n_12534;
or2_11085: n_12527 <=  n_12528  OR n_12531;
and2_11086: n_12528 <=  n_12529  AND n_12530;
inv_11087: n_12529  <= TRANSPORT NOT a_N2558_aNOT  ;
delay_11088: n_12530  <= TRANSPORT a_N2547  ;
and2_11089: n_12531 <=  n_12532  AND n_12533;
delay_11090: n_12532  <= TRANSPORT a_N2558_aNOT  ;
delay_11091: n_12533  <= TRANSPORT a_N183_aNOT  ;
and1_11092: n_12534 <=  gnd;
dff_11093: DFF_a8237

    PORT MAP ( D => a_EQ874, CLK => a_SCH0ADDRREG_F7_G_aCLK, CLRN => a_SCH0ADDRREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH0ADDRREG_F7_G);
inv_11094: a_SCH0ADDRREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11095: a_EQ874 <=  n_12541  XOR n_12552;
or3_11096: n_12541 <=  n_12542  OR n_12545  OR n_12548;
and2_11097: n_12542 <=  n_12543  AND n_12544;
inv_11098: n_12543  <= TRANSPORT NOT a_SCH0MODEREG_F2_G  ;
delay_11099: n_12544  <= TRANSPORT a_LC3_D9  ;
and2_11100: n_12545 <=  n_12546  AND n_12547;
inv_11101: n_12546  <= TRANSPORT NOT a_N57_aNOT  ;
delay_11102: n_12547  <= TRANSPORT a_LC3_D9  ;
and3_11103: n_12548 <=  n_12549  AND n_12550  AND n_12551;
delay_11104: n_12549  <= TRANSPORT a_N57_aNOT  ;
delay_11105: n_12550  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
delay_11106: n_12551  <= TRANSPORT a_SCH0BAROUT_F7_G  ;
and1_11107: n_12552 <=  gnd;
delay_11108: n_12553  <= TRANSPORT clk  ;
filter_11109: FILTER_a8237

    PORT MAP (IN1 => n_12553, Y => a_SCH0ADDRREG_F7_G_aCLK);
delay_11110: a_LC5_D19  <= TRANSPORT a_EQ685  ;
xor2_11111: a_EQ685 <=  n_12557  XOR n_12569;
or3_11112: n_12557 <=  n_12558  OR n_12562  OR n_12566;
and3_11113: n_12558 <=  n_12559  AND n_12560  AND n_12561;
inv_11114: n_12559  <= TRANSPORT NOT a_LC6_D6  ;
inv_11115: n_12560  <= TRANSPORT NOT a_N2352  ;
delay_11116: n_12561  <= TRANSPORT dbin(7)  ;
and2_11117: n_12562 <=  n_12563  AND n_12564;
delay_11118: n_12563  <= TRANSPORT a_N2352  ;
delay_11119: n_12564  <= TRANSPORT a_SCH1ADDRREG_F7_G  ;
and2_11120: n_12566 <=  n_12567  AND n_12568;
delay_11121: n_12567  <= TRANSPORT a_LC6_D6  ;
delay_11122: n_12568  <= TRANSPORT a_SCH1ADDRREG_F7_G  ;
and1_11123: n_12569 <=  gnd;
delay_11124: a_LC3_D19  <= TRANSPORT a_EQ686  ;
xor2_11125: a_EQ686 <=  n_12572  XOR n_12579;
or2_11126: n_12572 <=  n_12573  OR n_12576;
and2_11127: n_12573 <=  n_12574  AND n_12575;
inv_11128: n_12574  <= TRANSPORT NOT a_N2559_aNOT  ;
delay_11129: n_12575  <= TRANSPORT a_N2547  ;
and2_11130: n_12576 <=  n_12577  AND n_12578;
delay_11131: n_12577  <= TRANSPORT a_N2559_aNOT  ;
delay_11132: n_12578  <= TRANSPORT a_LC5_D19  ;
and1_11133: n_12579 <=  gnd;
dff_11134: DFF_a8237

    PORT MAP ( D => a_EQ938, CLK => a_SCH1ADDRREG_F7_G_aCLK, CLRN => a_SCH1ADDRREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCH1ADDRREG_F7_G);
inv_11135: a_SCH1ADDRREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11136: a_EQ938 <=  n_12586  XOR n_12597;
or3_11137: n_12586 <=  n_12587  OR n_12590  OR n_12593;
and2_11138: n_12587 <=  n_12588  AND n_12589;
inv_11139: n_12588  <= TRANSPORT NOT a_SCH1MODEREG_F2_G  ;
delay_11140: n_12589  <= TRANSPORT a_LC3_D19  ;
and2_11141: n_12590 <=  n_12591  AND n_12592;
inv_11142: n_12591  <= TRANSPORT NOT a_N57_aNOT  ;
delay_11143: n_12592  <= TRANSPORT a_LC3_D19  ;
and3_11144: n_12593 <=  n_12594  AND n_12595  AND n_12596;
delay_11145: n_12594  <= TRANSPORT a_N57_aNOT  ;
delay_11146: n_12595  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
delay_11147: n_12596  <= TRANSPORT a_SCH1BAROUT_F7_G  ;
and1_11148: n_12597 <=  gnd;
delay_11149: n_12598  <= TRANSPORT clk  ;
filter_11150: FILTER_a8237

    PORT MAP (IN1 => n_12598, Y => a_SCH1ADDRREG_F7_G_aCLK);
delay_11151: a_LC8_B25  <= TRANSPORT a_EQ430  ;
xor2_11152: a_EQ430 <=  n_12602  XOR n_12609;
or3_11153: n_12602 <=  n_12603  OR n_12605  OR n_12607;
and1_11154: n_12603 <=  n_12604;
delay_11155: n_12604  <= TRANSPORT a_N2372_aNOT  ;
and1_11156: n_12605 <=  n_12606;
delay_11157: n_12606  <= TRANSPORT a_N70  ;
and1_11158: n_12607 <=  n_12608;
inv_11159: n_12608  <= TRANSPORT NOT a_N2408_aNOT  ;
and1_11160: n_12609 <=  gnd;
delay_11161: a_N1467  <= TRANSPORT a_EQ448  ;
xor2_11162: a_EQ448 <=  n_12612  XOR n_12618;
or2_11163: n_12612 <=  n_12613  OR n_12616;
and2_11164: n_12613 <=  n_12614  AND n_12615;
inv_11165: n_12614  <= TRANSPORT NOT a_N822  ;
delay_11166: n_12615  <= TRANSPORT a_N821  ;
and1_11167: n_12616 <=  n_12617;
inv_11168: n_12617  <= TRANSPORT NOT a_N2374  ;
and1_11169: n_12618 <=  gnd;
dff_11170: DFF_a8237

    PORT MAP ( D => a_EQ306, CLK => a_N820_aCLK, CLRN => a_N820_aCLRN, PRN => vcc,
          Q => a_N820);
inv_11171: a_N820_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11172: a_EQ306 <=  n_12625  XOR n_12633;
or2_11173: n_12625 <=  n_12626  OR n_12629;
and2_11174: n_12626 <=  n_12627  AND n_12628;
delay_11175: n_12627  <= TRANSPORT a_N2563_aNOT  ;
delay_11176: n_12628  <= TRANSPORT a_LC8_B25  ;
and3_11177: n_12629 <=  n_12630  AND n_12631  AND n_12632;
delay_11178: n_12630  <= TRANSPORT a_N2563_aNOT  ;
delay_11179: n_12631  <= TRANSPORT a_N1467  ;
delay_11180: n_12632  <= TRANSPORT a_N820  ;
and1_11181: n_12633 <=  gnd;
delay_11182: n_12634  <= TRANSPORT clk  ;
filter_11183: FILTER_a8237

    PORT MAP (IN1 => n_12634, Y => a_N820_aCLK);
delay_11184: a_LC2_D4  <= TRANSPORT a_EQ360  ;
xor2_11185: a_EQ360 <=  n_12638  XOR n_12649;
or3_11186: n_12638 <=  n_12639  OR n_12642  OR n_12645;
and2_11187: n_12639 <=  n_12640  AND n_12641;
inv_11188: n_12640  <= TRANSPORT NOT a_LC3_E16_aNOT  ;
delay_11189: n_12641  <= TRANSPORT a_N3541  ;
and2_11190: n_12642 <=  n_12643  AND n_12644;
inv_11191: n_12643  <= TRANSPORT NOT a_N2557  ;
delay_11192: n_12644  <= TRANSPORT a_N3541  ;
and3_11193: n_12645 <=  n_12646  AND n_12647  AND n_12648;
delay_11194: n_12646  <= TRANSPORT a_N2557  ;
delay_11195: n_12647  <= TRANSPORT a_LC3_E16_aNOT  ;
inv_11196: n_12648  <= TRANSPORT NOT a_N3541  ;
and1_11197: n_12649 <=  gnd;
delay_11198: a_N1141  <= TRANSPORT a_EQ367  ;
xor2_11199: a_EQ367 <=  n_12652  XOR n_12659;
or2_11200: n_12652 <=  n_12653  OR n_12656;
and2_11201: n_12653 <=  n_12654  AND n_12655;
delay_11202: n_12654  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_11203: n_12655  <= TRANSPORT a_SH1WRDCNTREG_F15_G  ;
and2_11204: n_12656 <=  n_12657  AND n_12658;
inv_11205: n_12657  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_11206: n_12658  <= TRANSPORT a_SH0WRDCNTREG_F15_G  ;
and1_11207: n_12659 <=  gnd;
delay_11208: a_LC1_D4  <= TRANSPORT a_EQ366  ;
xor2_11209: a_EQ366 <=  n_12662  XOR n_12669;
or2_11210: n_12662 <=  n_12663  OR n_12666;
and2_11211: n_12663 <=  n_12664  AND n_12665;
inv_11212: n_12664  <= TRANSPORT NOT a_N2531  ;
delay_11213: n_12665  <= TRANSPORT a_LC2_D4  ;
and2_11214: n_12666 <=  n_12667  AND n_12668;
delay_11215: n_12667  <= TRANSPORT a_N2531  ;
delay_11216: n_12668  <= TRANSPORT a_N1141  ;
and1_11217: n_12669 <=  gnd;
delay_11218: a_LC4_D12  <= TRANSPORT a_EQ369  ;
xor2_11219: a_EQ369 <=  n_12672  XOR n_12679;
or2_11220: n_12672 <=  n_12673  OR n_12676;
and2_11221: n_12673 <=  n_12674  AND n_12675;
inv_11222: n_12674  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_11223: n_12675  <= TRANSPORT a_SH0WRDCNTREG_F15_G  ;
and2_11224: n_12676 <=  n_12677  AND n_12678;
inv_11225: n_12677  <= TRANSPORT NOT a_N88_aNOT  ;
delay_11226: n_12678  <= TRANSPORT a_SH1WRDCNTREG_F15_G  ;
and1_11227: n_12679 <=  gnd;
delay_11228: a_LC3_D12  <= TRANSPORT a_EQ368  ;
xor2_11229: a_EQ368 <=  n_12682  XOR n_12689;
or2_11230: n_12682 <=  n_12683  OR n_12686;
and2_11231: n_12683 <=  n_12684  AND n_12685;
inv_11232: n_12684  <= TRANSPORT NOT a_N2376  ;
delay_11233: n_12685  <= TRANSPORT a_SH2WRDCNTREG_F15_G  ;
and2_11234: n_12686 <=  n_12687  AND n_12688;
inv_11235: n_12687  <= TRANSPORT NOT a_N2377  ;
delay_11236: n_12688  <= TRANSPORT a_SH3WRDCNTREG_F15_G  ;
and1_11237: n_12689 <=  gnd;
dff_11238: DFF_a8237

    PORT MAP ( D => a_EQ837, CLK => a_N3541_aCLK, CLRN => a_N3541_aCLRN, PRN => vcc,
          Q => a_N3541);
inv_11239: a_N3541_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11240: a_EQ837 <=  n_12696  XOR n_12706;
or3_11241: n_12696 <=  n_12697  OR n_12700  OR n_12703;
and2_11242: n_12697 <=  n_12698  AND n_12699;
delay_11243: n_12698  <= TRANSPORT a_LC1_D4  ;
inv_11244: n_12699  <= TRANSPORT NOT startdma  ;
and2_11245: n_12700 <=  n_12701  AND n_12702;
delay_11246: n_12701  <= TRANSPORT a_LC4_D12  ;
delay_11247: n_12702  <= TRANSPORT startdma  ;
and2_11248: n_12703 <=  n_12704  AND n_12705;
delay_11249: n_12704  <= TRANSPORT a_LC3_D12  ;
delay_11250: n_12705  <= TRANSPORT startdma  ;
and1_11251: n_12706 <=  gnd;
delay_11252: n_12707  <= TRANSPORT clk  ;
filter_11253: FILTER_a8237

    PORT MAP (IN1 => n_12707, Y => a_N3541_aCLK);
delay_11254: a_N2395  <= TRANSPORT a_N2395_aIN  ;
xor2_11255: a_N2395_aIN <=  n_12711  XOR n_12716;
or1_11256: n_12711 <=  n_12712;
and3_11257: n_12712 <=  n_12713  AND n_12714  AND n_12715;
inv_11258: n_12713  <= TRANSPORT NOT a_N71_aNOT  ;
inv_11259: n_12714  <= TRANSPORT NOT a_N2539  ;
inv_11260: n_12715  <= TRANSPORT NOT a_N825  ;
and1_11261: n_12716 <=  gnd;
delay_11262: a_LC4_B13  <= TRANSPORT a_EQ392  ;
xor2_11263: a_EQ392 <=  n_12719  XOR n_12726;
or3_11264: n_12719 <=  n_12720  OR n_12722  OR n_12724;
and1_11265: n_12720 <=  n_12721;
delay_11266: n_12721  <= TRANSPORT a_N70  ;
and1_11267: n_12722 <=  n_12723;
inv_11268: n_12723  <= TRANSPORT NOT a_N2358  ;
and1_11269: n_12724 <=  n_12725;
delay_11270: n_12725  <= TRANSPORT a_N2395  ;
and1_11271: n_12726 <=  gnd;
dff_11272: DFF_a8237

    PORT MAP ( D => a_N4179_aD, CLK => a_N4179_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4179);
xor2_11273: a_N4179_aD <=  n_12734  XOR n_12737;
or1_11274: n_12734 <=  n_12735;
and1_11275: n_12735 <=  n_12736;
delay_11276: n_12736  <= TRANSPORT dreq(2)  ;
and1_11277: n_12737 <=  gnd;
delay_11278: n_12738  <= TRANSPORT clk  ;
filter_11279: FILTER_a8237

    PORT MAP (IN1 => n_12738, Y => a_N4179_aCLK);
dff_11280: DFF_a8237

    PORT MAP ( D => a_N4183_aD, CLK => a_N4183_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4183);
xor2_11281: a_N4183_aD <=  n_12746  XOR n_12749;
or1_11282: n_12746 <=  n_12747;
and1_11283: n_12747 <=  n_12748;
delay_11284: n_12748  <= TRANSPORT a_N4179  ;
and1_11285: n_12749 <=  gnd;
delay_11286: n_12750  <= TRANSPORT clk  ;
filter_11287: FILTER_a8237

    PORT MAP (IN1 => n_12750, Y => a_N4183_aCLK);
delay_11288: a_N59  <= TRANSPORT a_EQ182  ;
xor2_11289: a_EQ182 <=  n_12754  XOR n_12766;
or3_11290: n_12754 <=  n_12755  OR n_12759  OR n_12763;
and3_11291: n_12755 <=  n_12756  AND n_12757  AND n_12758;
inv_11292: n_12756  <= TRANSPORT NOT a_SREQUESTREG_F2_G  ;
inv_11293: n_12757  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
inv_11294: n_12758  <= TRANSPORT NOT a_N4183  ;
and3_11295: n_12759 <=  n_12760  AND n_12761  AND n_12762;
inv_11296: n_12760  <= TRANSPORT NOT a_SREQUESTREG_F2_G  ;
delay_11297: n_12761  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
delay_11298: n_12762  <= TRANSPORT a_N4183  ;
and2_11299: n_12763 <=  n_12764  AND n_12765;
inv_11300: n_12764  <= TRANSPORT NOT a_SREQUESTREG_F2_G  ;
inv_11301: n_12765  <= TRANSPORT NOT a_SMASKREG_F2_G_aNOT  ;
and1_11302: n_12766 <=  gnd;
dff_11303: DFF_a8237

    PORT MAP ( D => a_N4178_aD, CLK => a_N4178_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4178);
xor2_11304: a_N4178_aD <=  n_12774  XOR n_12777;
or1_11305: n_12774 <=  n_12775;
and1_11306: n_12775 <=  n_12776;
delay_11307: n_12776  <= TRANSPORT dreq(3)  ;
and1_11308: n_12777 <=  gnd;
delay_11309: n_12778  <= TRANSPORT clk  ;
filter_11310: FILTER_a8237

    PORT MAP (IN1 => n_12778, Y => a_N4178_aCLK);
dff_11311: DFF_a8237

    PORT MAP ( D => a_N4182_aD, CLK => a_N4182_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4182);
xor2_11312: a_N4182_aD <=  n_12786  XOR n_12789;
or1_11313: n_12786 <=  n_12787;
and1_11314: n_12787 <=  n_12788;
delay_11315: n_12788  <= TRANSPORT a_N4178  ;
and1_11316: n_12789 <=  gnd;
delay_11317: n_12790  <= TRANSPORT clk  ;
filter_11318: FILTER_a8237

    PORT MAP (IN1 => n_12790, Y => a_N4182_aCLK);
delay_11319: a_N2534  <= TRANSPORT a_EQ594  ;
xor2_11320: a_EQ594 <=  n_12794  XOR n_12805;
or3_11321: n_12794 <=  n_12795  OR n_12799  OR n_12803;
and3_11322: n_12795 <=  n_12796  AND n_12797  AND n_12798;
delay_11323: n_12796  <= TRANSPORT a_SMASKREG_F3_G_aNOT  ;
inv_11324: n_12797  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
delay_11325: n_12798  <= TRANSPORT a_N4182  ;
and3_11326: n_12799 <=  n_12800  AND n_12801  AND n_12802;
delay_11327: n_12800  <= TRANSPORT a_SMASKREG_F3_G_aNOT  ;
delay_11328: n_12801  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
inv_11329: n_12802  <= TRANSPORT NOT a_N4182  ;
and1_11330: n_12803 <=  n_12804;
delay_11331: n_12804  <= TRANSPORT a_SREQUESTREG_F3_G  ;
and1_11332: n_12805 <=  gnd;
delay_11333: a_LC3_B6  <= TRANSPORT a_EQ596  ;
xor2_11334: a_EQ596 <=  n_12808  XOR n_12815;
or2_11335: n_12808 <=  n_12809  OR n_12812;
and2_11336: n_12809 <=  n_12810  AND n_12811;
inv_11337: n_12810  <= TRANSPORT NOT a_N2376  ;
inv_11338: n_12811  <= TRANSPORT NOT a_N59  ;
and2_11339: n_12812 <=  n_12813  AND n_12814;
inv_11340: n_12813  <= TRANSPORT NOT a_N2377  ;
delay_11341: n_12814  <= TRANSPORT a_N2534  ;
and1_11342: n_12815 <=  gnd;
delay_11343: a_LC4_E2  <= TRANSPORT a_EQ474  ;
xor2_11344: a_EQ474 <=  n_12818  XOR n_12831;
or4_11345: n_12818 <=  n_12819  OR n_12822  OR n_12825  OR n_12828;
and2_11346: n_12819 <=  n_12820  AND n_12821;
inv_11347: n_12820  <= TRANSPORT NOT a_SCH2MODEREG_F4_G  ;
inv_11348: n_12821  <= TRANSPORT NOT a_SCH3MODEREG_F4_G  ;
and2_11349: n_12822 <=  n_12823  AND n_12824;
delay_11350: n_12823  <= TRANSPORT a_N2377  ;
inv_11351: n_12824  <= TRANSPORT NOT a_SCH2MODEREG_F4_G  ;
and2_11352: n_12825 <=  n_12826  AND n_12827;
delay_11353: n_12826  <= TRANSPORT a_N2376  ;
inv_11354: n_12827  <= TRANSPORT NOT a_SCH3MODEREG_F4_G  ;
and2_11355: n_12828 <=  n_12829  AND n_12830;
delay_11356: n_12829  <= TRANSPORT a_N2377  ;
delay_11357: n_12830  <= TRANSPORT a_N2376  ;
and1_11358: n_12831 <=  gnd;
delay_11359: a_LC1_E2  <= TRANSPORT a_EQ473  ;
xor2_11360: a_EQ473 <=  n_12834  XOR n_12847;
or4_11361: n_12834 <=  n_12835  OR n_12838  OR n_12841  OR n_12844;
and2_11362: n_12835 <=  n_12836  AND n_12837;
inv_11363: n_12836  <= TRANSPORT NOT a_SCH1MODEREG_F4_G  ;
inv_11364: n_12837  <= TRANSPORT NOT a_SCH0MODEREG_F4_G  ;
and2_11365: n_12838 <=  n_12839  AND n_12840;
delay_11366: n_12839  <= TRANSPORT a_N88_aNOT  ;
inv_11367: n_12840  <= TRANSPORT NOT a_SCH0MODEREG_F4_G  ;
and2_11368: n_12841 <=  n_12842  AND n_12843;
delay_11369: n_12842  <= TRANSPORT a_N2598_aNOT  ;
inv_11370: n_12843  <= TRANSPORT NOT a_SCH1MODEREG_F4_G  ;
and2_11371: n_12844 <=  n_12845  AND n_12846;
delay_11372: n_12845  <= TRANSPORT a_N2598_aNOT  ;
delay_11373: n_12846  <= TRANSPORT a_N88_aNOT  ;
and1_11374: n_12847 <=  gnd;
dff_11375: DFF_a8237

    PORT MAP ( D => a_N4180_aD, CLK => a_N4180_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4180);
xor2_11376: a_N4180_aD <=  n_12855  XOR n_12858;
or1_11377: n_12855 <=  n_12856;
and1_11378: n_12856 <=  n_12857;
delay_11379: n_12857  <= TRANSPORT dreq(1)  ;
and1_11380: n_12858 <=  gnd;
delay_11381: n_12859  <= TRANSPORT clk  ;
filter_11382: FILTER_a8237

    PORT MAP (IN1 => n_12859, Y => a_N4180_aCLK);
dff_11383: DFF_a8237

    PORT MAP ( D => a_N4184_aD, CLK => a_N4184_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4184);
xor2_11384: a_N4184_aD <=  n_12867  XOR n_12870;
or1_11385: n_12867 <=  n_12868;
and1_11386: n_12868 <=  n_12869;
delay_11387: n_12869  <= TRANSPORT a_N4180  ;
and1_11388: n_12870 <=  gnd;
delay_11389: n_12871  <= TRANSPORT clk  ;
filter_11390: FILTER_a8237

    PORT MAP (IN1 => n_12871, Y => a_N4184_aCLK);
delay_11391: a_N2536  <= TRANSPORT a_EQ595  ;
xor2_11392: a_EQ595 <=  n_12875  XOR n_12886;
or3_11393: n_12875 <=  n_12876  OR n_12880  OR n_12884;
and3_11394: n_12876 <=  n_12877  AND n_12878  AND n_12879;
delay_11395: n_12877  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
delay_11396: n_12878  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
inv_11397: n_12879  <= TRANSPORT NOT a_N4184  ;
and3_11398: n_12880 <=  n_12881  AND n_12882  AND n_12883;
delay_11399: n_12881  <= TRANSPORT a_SMASKREG_F1_G_aNOT  ;
inv_11400: n_12882  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
delay_11401: n_12883  <= TRANSPORT a_N4184  ;
and1_11402: n_12884 <=  n_12885;
delay_11403: n_12885  <= TRANSPORT a_SREQUESTREG_F1_G  ;
and1_11404: n_12886 <=  gnd;
dff_11405: DFF_a8237

    PORT MAP ( D => a_N4181_aD, CLK => a_N4181_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4181);
xor2_11406: a_N4181_aD <=  n_12894  XOR n_12897;
or1_11407: n_12894 <=  n_12895;
and1_11408: n_12895 <=  n_12896;
delay_11409: n_12896  <= TRANSPORT dreq(0)  ;
and1_11410: n_12897 <=  gnd;
delay_11411: n_12898  <= TRANSPORT clk  ;
filter_11412: FILTER_a8237

    PORT MAP (IN1 => n_12898, Y => a_N4181_aCLK);
dff_11413: DFF_a8237

    PORT MAP ( D => a_N4185_aD, CLK => a_N4185_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4185);
xor2_11414: a_N4185_aD <=  n_12906  XOR n_12909;
or1_11415: n_12906 <=  n_12907;
and1_11416: n_12907 <=  n_12908;
delay_11417: n_12908  <= TRANSPORT a_N4181  ;
and1_11418: n_12909 <=  gnd;
delay_11419: n_12910  <= TRANSPORT clk  ;
filter_11420: FILTER_a8237

    PORT MAP (IN1 => n_12910, Y => a_N4185_aCLK);
delay_11421: a_N55  <= TRANSPORT a_EQ180  ;
xor2_11422: a_EQ180 <=  n_12914  XOR n_12926;
or3_11423: n_12914 <=  n_12915  OR n_12919  OR n_12923;
and3_11424: n_12915 <=  n_12916  AND n_12917  AND n_12918;
inv_11425: n_12916  <= TRANSPORT NOT a_SREQUESTREG_F0_G  ;
delay_11426: n_12917  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
delay_11427: n_12918  <= TRANSPORT a_N4185  ;
and3_11428: n_12919 <=  n_12920  AND n_12921  AND n_12922;
inv_11429: n_12920  <= TRANSPORT NOT a_SREQUESTREG_F0_G  ;
inv_11430: n_12921  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
inv_11431: n_12922  <= TRANSPORT NOT a_N4185  ;
and2_11432: n_12923 <=  n_12924  AND n_12925;
inv_11433: n_12924  <= TRANSPORT NOT a_SMASKREG_F0_G_aNOT  ;
inv_11434: n_12925  <= TRANSPORT NOT a_SREQUESTREG_F0_G  ;
and1_11435: n_12926 <=  gnd;
delay_11436: a_LC4_B16  <= TRANSPORT a_EQ597  ;
xor2_11437: a_EQ597 <=  n_12929  XOR n_12936;
or2_11438: n_12929 <=  n_12930  OR n_12933;
and2_11439: n_12930 <=  n_12931  AND n_12932;
inv_11440: n_12931  <= TRANSPORT NOT a_N88_aNOT  ;
delay_11441: n_12932  <= TRANSPORT a_N2536  ;
and2_11442: n_12933 <=  n_12934  AND n_12935;
inv_11443: n_12934  <= TRANSPORT NOT a_N2598_aNOT  ;
inv_11444: n_12935  <= TRANSPORT NOT a_N55  ;
and1_11445: n_12936 <=  gnd;
delay_11446: a_N1585_aNOT  <= TRANSPORT a_EQ475  ;
xor2_11447: a_EQ475 <=  n_12939  XOR n_12948;
or2_11448: n_12939 <=  n_12940  OR n_12944;
and3_11449: n_12940 <=  n_12941  AND n_12942  AND n_12943;
delay_11450: n_12941  <= TRANSPORT a_LC3_B6  ;
delay_11451: n_12942  <= TRANSPORT a_LC4_E2  ;
delay_11452: n_12943  <= TRANSPORT a_LC1_E2  ;
and3_11453: n_12944 <=  n_12945  AND n_12946  AND n_12947;
delay_11454: n_12945  <= TRANSPORT a_LC4_E2  ;
delay_11455: n_12946  <= TRANSPORT a_LC1_E2  ;
delay_11456: n_12947  <= TRANSPORT a_LC4_B16  ;
and1_11457: n_12948 <=  gnd;
delay_11458: a_LC1_E15  <= TRANSPORT a_EQ469  ;
xor2_11459: a_EQ469 <=  n_12951  XOR n_12958;
or2_11460: n_12951 <=  n_12952  OR n_12955;
and2_11461: n_12952 <=  n_12953  AND n_12954;
inv_11462: n_12953  <= TRANSPORT NOT a_N88_aNOT  ;
delay_11463: n_12954  <= TRANSPORT a_SCH1MODEREG_F5_G  ;
and2_11464: n_12955 <=  n_12956  AND n_12957;
inv_11465: n_12956  <= TRANSPORT NOT a_N2377  ;
delay_11466: n_12957  <= TRANSPORT a_SCH3MODEREG_F5_G  ;
and1_11467: n_12958 <=  gnd;
delay_11468: a_LC6_E26  <= TRANSPORT a_EQ470  ;
xor2_11469: a_EQ470 <=  n_12961  XOR n_12968;
or2_11470: n_12961 <=  n_12962  OR n_12965;
and2_11471: n_12962 <=  n_12963  AND n_12964;
inv_11472: n_12963  <= TRANSPORT NOT a_N2376  ;
delay_11473: n_12964  <= TRANSPORT a_SCH2MODEREG_F5_G  ;
and2_11474: n_12965 <=  n_12966  AND n_12967;
inv_11475: n_12966  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_11476: n_12967  <= TRANSPORT a_SCH0MODEREG_F5_G  ;
and1_11477: n_12968 <=  gnd;
delay_11478: a_N1581_aNOT  <= TRANSPORT a_EQ471  ;
xor2_11479: a_EQ471 <=  n_12971  XOR n_12978;
or3_11480: n_12971 <=  n_12972  OR n_12974  OR n_12976;
and1_11481: n_12972 <=  n_12973;
delay_11482: n_12973  <= TRANSPORT a_N1585_aNOT  ;
and1_11483: n_12974 <=  n_12975;
delay_11484: n_12975  <= TRANSPORT a_LC1_E15  ;
and1_11485: n_12976 <=  n_12977;
delay_11486: n_12977  <= TRANSPORT a_LC6_E26  ;
and1_11487: n_12978 <=  gnd;
delay_11488: a_N2394  <= TRANSPORT a_N2394_aIN  ;
xor2_11489: a_N2394_aIN <=  n_12981  XOR n_12987;
or1_11490: n_12981 <=  n_12982;
and4_11491: n_12982 <=  n_12983  AND n_12984  AND n_12985  AND n_12986;
inv_11492: n_12983  <= TRANSPORT NOT a_N2361  ;
inv_11493: n_12984  <= TRANSPORT NOT a_N2539  ;
inv_11494: n_12985  <= TRANSPORT NOT a_N825  ;
delay_11495: n_12986  <= TRANSPORT a_N1581_aNOT  ;
and1_11496: n_12987 <=  gnd;
delay_11497: a_N2369_aNOT  <= TRANSPORT a_N2369_aNOT_aIN  ;
xor2_11498: a_N2369_aNOT_aIN <=  n_12990  XOR n_12996;
or1_11499: n_12990 <=  n_12991;
and4_11500: n_12991 <=  n_12992  AND n_12993  AND n_12994  AND n_12995;
inv_11501: n_12992  <= TRANSPORT NOT a_LC4_E22  ;
delay_11502: n_12993  <= TRANSPORT a_LC6_E22  ;
delay_11503: n_12994  <= TRANSPORT a_LC5_E22  ;
inv_11504: n_12995  <= TRANSPORT NOT a_LC6_E10  ;
and1_11505: n_12996 <=  gnd;
delay_11506: a_LC4_B3  <= TRANSPORT a_EQ393  ;
xor2_11507: a_EQ393 <=  n_13000  XOR n_13010;
or3_11508: n_13000 <=  n_13001  OR n_13004  OR n_13007;
and2_11509: n_13001 <=  n_13002  AND n_13003;
inv_11510: n_13002  <= TRANSPORT NOT a_N2356  ;
delay_11511: n_13003  <= TRANSPORT a_N2369_aNOT  ;
and2_11512: n_13004 <=  n_13005  AND n_13006;
inv_11513: n_13005  <= TRANSPORT NOT a_N2356  ;
delay_11514: n_13006  <= TRANSPORT ready  ;
and2_11515: n_13007 <=  n_13008  AND n_13009;
inv_11516: n_13008  <= TRANSPORT NOT a_N67_aNOT  ;
delay_11517: n_13009  <= TRANSPORT ready  ;
and1_11518: n_13010 <=  gnd;
delay_11519: a_N2359_aNOT  <= TRANSPORT a_N2359_aNOT_aIN  ;
xor2_11520: a_N2359_aNOT_aIN <=  n_13013  XOR n_13017;
or1_11521: n_13013 <=  n_13014;
and2_11522: n_13014 <=  n_13015  AND n_13016;
inv_11523: n_13015  <= TRANSPORT NOT a_N1566  ;
delay_11524: n_13016  <= TRANSPORT a_N823  ;
and1_11525: n_13017 <=  gnd;
delay_11526: a_LC3_B16  <= TRANSPORT a_EQ394  ;
xor2_11527: a_EQ394 <=  n_13020  XOR n_13027;
or2_11528: n_13020 <=  n_13021  OR n_13024;
and2_11529: n_13021 <=  n_13022  AND n_13023;
inv_11530: n_13022  <= TRANSPORT NOT a_N68_aNOT  ;
delay_11531: n_13023  <= TRANSPORT a_SCOMMANDREG_F3_G  ;
and2_11532: n_13024 <=  n_13025  AND n_13026;
delay_11533: n_13025  <= TRANSPORT a_N2359_aNOT  ;
delay_11534: n_13026  <= TRANSPORT startdma  ;
and1_11535: n_13027 <=  gnd;
delay_11536: a_N1249  <= TRANSPORT a_N1249_aIN  ;
xor2_11537: a_N1249_aIN <=  n_13030  XOR n_13036;
or1_11538: n_13030 <=  n_13031;
and4_11539: n_13031 <=  n_13032  AND n_13033  AND n_13034  AND n_13035;
delay_11540: n_13032  <= TRANSPORT a_N820  ;
inv_11541: n_13033  <= TRANSPORT NOT a_N822  ;
delay_11542: n_13034  <= TRANSPORT a_N821  ;
delay_11543: n_13035  <= TRANSPORT a_N823  ;
and1_11544: n_13036 <=  gnd;
delay_11545: a_LC3_B3  <= TRANSPORT a_EQ395  ;
xor2_11546: a_EQ395 <=  n_13039  XOR n_13048;
or4_11547: n_13039 <=  n_13040  OR n_13042  OR n_13044  OR n_13046;
and1_11548: n_13040 <=  n_13041;
delay_11549: n_13041  <= TRANSPORT a_LC4_B3  ;
and1_11550: n_13042 <=  n_13043;
delay_11551: n_13043  <= TRANSPORT a_LC3_B16  ;
and1_11552: n_13044 <=  n_13045;
delay_11553: n_13045  <= TRANSPORT a_N1249  ;
and1_11554: n_13046 <=  n_13047;
delay_11555: n_13047  <= TRANSPORT a_N2372_aNOT  ;
and1_11556: n_13048 <=  gnd;
dff_11557: DFF_a8237

    PORT MAP ( D => a_EQ308, CLK => a_N822_aCLK, CLRN => a_N822_aCLRN, PRN => vcc,
          Q => a_N822);
inv_11558: a_N822_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11559: a_EQ308 <=  n_13055  XOR n_13065;
or3_11560: n_13055 <=  n_13056  OR n_13059  OR n_13062;
and2_11561: n_13056 <=  n_13057  AND n_13058;
delay_11562: n_13057  <= TRANSPORT a_N2563_aNOT  ;
delay_11563: n_13058  <= TRANSPORT a_LC4_B13  ;
and2_11564: n_13059 <=  n_13060  AND n_13061;
delay_11565: n_13060  <= TRANSPORT a_N2563_aNOT  ;
delay_11566: n_13061  <= TRANSPORT a_N2394  ;
and2_11567: n_13062 <=  n_13063  AND n_13064;
delay_11568: n_13063  <= TRANSPORT a_N2563_aNOT  ;
delay_11569: n_13064  <= TRANSPORT a_LC3_B3  ;
and1_11570: n_13065 <=  gnd;
delay_11571: n_13066  <= TRANSPORT clk  ;
filter_11572: FILTER_a8237

    PORT MAP (IN1 => n_13066, Y => a_N822_aCLK);
delay_11573: a_N1387  <= TRANSPORT a_N1387_aIN  ;
xor2_11574: a_N1387_aIN <=  n_13070  XOR n_13075;
or1_11575: n_13070 <=  n_13071;
and3_11576: n_13071 <=  n_13072  AND n_13073  AND n_13074;
delay_11577: n_13072  <= TRANSPORT a_N2591  ;
delay_11578: n_13073  <= TRANSPORT a_N2359_aNOT  ;
delay_11579: n_13074  <= TRANSPORT startdma  ;
and1_11580: n_13075 <=  gnd;
delay_11581: a_LC8_B13  <= TRANSPORT a_EQ429  ;
xor2_11582: a_EQ429 <=  n_13078  XOR n_13086;
or2_11583: n_13078 <=  n_13079  OR n_13082;
and2_11584: n_13079 <=  n_13080  AND n_13081;
inv_11585: n_13080  <= TRANSPORT NOT a_N822  ;
delay_11586: n_13081  <= TRANSPORT a_N821  ;
and3_11587: n_13082 <=  n_13083  AND n_13084  AND n_13085;
delay_11588: n_13083  <= TRANSPORT a_N822  ;
inv_11589: n_13084  <= TRANSPORT NOT a_N821  ;
delay_11590: n_13085  <= TRANSPORT a_N823  ;
and1_11591: n_13086 <=  gnd;
dff_11592: DFF_a8237

    PORT MAP ( D => a_EQ307, CLK => a_N821_aCLK, CLRN => a_N821_aCLRN, PRN => vcc,
          Q => a_N821);
inv_11593: a_N821_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11594: a_EQ307 <=  n_13093  XOR n_13103;
or3_11595: n_13093 <=  n_13094  OR n_13097  OR n_13100;
and2_11596: n_13094 <=  n_13095  AND n_13096;
delay_11597: n_13095  <= TRANSPORT a_N2563_aNOT  ;
delay_11598: n_13096  <= TRANSPORT a_N2395  ;
and2_11599: n_13097 <=  n_13098  AND n_13099;
delay_11600: n_13098  <= TRANSPORT a_N2563_aNOT  ;
delay_11601: n_13099  <= TRANSPORT a_N1387  ;
and2_11602: n_13100 <=  n_13101  AND n_13102;
delay_11603: n_13101  <= TRANSPORT a_N2563_aNOT  ;
delay_11604: n_13102  <= TRANSPORT a_LC8_B13  ;
and1_11605: n_13103 <=  gnd;
delay_11606: n_13104  <= TRANSPORT clk  ;
filter_11607: FILTER_a8237

    PORT MAP (IN1 => n_13104, Y => a_N821_aCLK);
dff_11608: DFF_a8237

    PORT MAP ( D => a_EQ1185, CLK => a_STEMPORARYREG_F4_G_aCLK, CLRN => a_STEMPORARYREG_F4_G_aCLRN,
          PRN => vcc, Q => a_STEMPORARYREG_F4_G);
inv_11609: a_STEMPORARYREG_F4_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11610: a_EQ1185 <=  n_13113  XOR n_13122;
or2_11611: n_13113 <=  n_13114  OR n_13118;
and3_11612: n_13114 <=  n_13115  AND n_13116  AND n_13117;
delay_11613: n_13115  <= TRANSPORT a_N2563_aNOT  ;
inv_11614: n_13116  <= TRANSPORT NOT a_N2372_aNOT  ;
delay_11615: n_13117  <= TRANSPORT a_STEMPORARYREG_F4_G  ;
and3_11616: n_13118 <=  n_13119  AND n_13120  AND n_13121;
delay_11617: n_13119  <= TRANSPORT a_N2563_aNOT  ;
delay_11618: n_13120  <= TRANSPORT a_N2372_aNOT  ;
delay_11619: n_13121  <= TRANSPORT dbin(4)  ;
and1_11620: n_13122 <=  gnd;
delay_11621: n_13123  <= TRANSPORT clk  ;
filter_11622: FILTER_a8237

    PORT MAP (IN1 => n_13123, Y => a_STEMPORARYREG_F4_G_aCLK);
dff_11623: DFF_a8237

    PORT MAP ( D => a_EQ1130, CLK => a_SCOMMANDREG_F7_G_aCLK, CLRN => a_SCOMMANDREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F7_G);
inv_11624: a_SCOMMANDREG_F7_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11625: a_EQ1130 <=  n_13132  XOR n_13141;
or2_11626: n_13132 <=  n_13133  OR n_13137;
and3_11627: n_13133 <=  n_13134  AND n_13135  AND n_13136;
delay_11628: n_13134  <= TRANSPORT a_N2563_aNOT  ;
delay_11629: n_13135  <= TRANSPORT a_N2571_aNOT  ;
delay_11630: n_13136  <= TRANSPORT a_SCOMMANDREG_F7_G  ;
and3_11631: n_13137 <=  n_13138  AND n_13139  AND n_13140;
delay_11632: n_13138  <= TRANSPORT a_N2563_aNOT  ;
inv_11633: n_13139  <= TRANSPORT NOT a_N2571_aNOT  ;
delay_11634: n_13140  <= TRANSPORT dbin(7)  ;
and1_11635: n_13141 <=  gnd;
delay_11636: n_13142  <= TRANSPORT clk  ;
filter_11637: FILTER_a8237

    PORT MAP (IN1 => n_13142, Y => a_SCOMMANDREG_F7_G_aCLK);
delay_11638: a_N2606  <= TRANSPORT a_EQ648  ;
xor2_11639: a_EQ648 <=  n_13146  XOR n_13151;
or2_11640: n_13146 <=  n_13147  OR n_13149;
and1_11641: n_13147 <=  n_13148;
inv_11642: n_13148  <= TRANSPORT NOT a_N59  ;
and1_11643: n_13149 <=  n_13150;
delay_11644: n_13150  <= TRANSPORT a_N2534  ;
and1_11645: n_13151 <=  gnd;
delay_11646: a_LC2_B2  <= TRANSPORT a_EQ543  ;
xor2_11647: a_EQ543 <=  n_13154  XOR n_13162;
or2_11648: n_13154 <=  n_13155  OR n_13159;
and3_11649: n_13155 <=  n_13156  AND n_13157  AND n_13158;
inv_11650: n_13156  <= TRANSPORT NOT a_N2598_aNOT  ;
inv_11651: n_13157  <= TRANSPORT NOT a_N2536  ;
delay_11652: n_13158  <= TRANSPORT a_N2606  ;
and2_11653: n_13159 <=  n_13160  AND n_13161;
inv_11654: n_13160  <= TRANSPORT NOT a_N88_aNOT  ;
delay_11655: n_13161  <= TRANSPORT a_N2606  ;
and1_11656: n_13162 <=  gnd;
delay_11657: a_LC6_B2  <= TRANSPORT a_EQ544  ;
xor2_11658: a_EQ544 <=  n_13165  XOR n_13172;
or2_11659: n_13165 <=  n_13166  OR n_13170;
and3_11660: n_13166 <=  n_13167  AND n_13168  AND n_13169;
inv_11661: n_13167  <= TRANSPORT NOT a_N59  ;
inv_11662: n_13168  <= TRANSPORT NOT a_N2536  ;
delay_11663: n_13169  <= TRANSPORT a_N55  ;
and1_11664: n_13170 <=  n_13171;
delay_11665: n_13171  <= TRANSPORT a_N2534  ;
and1_11666: n_13172 <=  gnd;
delay_11667: a_LC7_B2  <= TRANSPORT a_EQ545  ;
xor2_11668: a_EQ545 <=  n_13175  XOR n_13183;
or2_11669: n_13175 <=  n_13176  OR n_13179;
and2_11670: n_13176 <=  n_13177  AND n_13178;
delay_11671: n_13177  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
delay_11672: n_13178  <= TRANSPORT a_LC2_B2  ;
and3_11673: n_13179 <=  n_13180  AND n_13181  AND n_13182;
inv_11674: n_13180  <= TRANSPORT NOT a_N2376  ;
delay_11675: n_13181  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
delay_11676: n_13182  <= TRANSPORT a_LC6_B2  ;
and1_11677: n_13183 <=  gnd;
delay_11678: a_LC5_B2  <= TRANSPORT a_EQ542  ;
xor2_11679: a_EQ542 <=  n_13186  XOR n_13193;
or2_11680: n_13186 <=  n_13187  OR n_13190;
and2_11681: n_13187 <=  n_13188  AND n_13189;
inv_11682: n_13188  <= TRANSPORT NOT a_SCOMMANDREG_F4_G  ;
delay_11683: n_13189  <= TRANSPORT a_N2606  ;
and2_11684: n_13190 <=  n_13191  AND n_13192;
inv_11685: n_13191  <= TRANSPORT NOT a_N2377  ;
delay_11686: n_13192  <= TRANSPORT a_N2606  ;
and1_11687: n_13193 <=  gnd;
delay_11688: a_LC4_B2  <= TRANSPORT a_EQ546  ;
xor2_11689: a_EQ546 <=  n_13196  XOR n_13203;
or2_11690: n_13196 <=  n_13197  OR n_13199;
and1_11691: n_13197 <=  n_13198;
delay_11692: n_13198  <= TRANSPORT a_LC7_B2  ;
and3_11693: n_13199 <=  n_13200  AND n_13201  AND n_13202;
inv_11694: n_13200  <= TRANSPORT NOT a_N2536  ;
delay_11695: n_13201  <= TRANSPORT a_N55  ;
delay_11696: n_13202  <= TRANSPORT a_LC5_B2  ;
and1_11697: n_13203 <=  gnd;
dff_11698: DFF_a8237

    PORT MAP ( D => a_N4186_aD, CLK => a_N4186_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4186);
xor2_11699: a_N4186_aD <=  n_13211  XOR n_13214;
or1_11700: n_13211 <=  n_13212;
and1_11701: n_13212 <=  n_13213;
delay_11702: n_13213  <= TRANSPORT hlda  ;
and1_11703: n_13214 <=  gnd;
delay_11704: n_13215  <= TRANSPORT clk  ;
filter_11705: FILTER_a8237

    PORT MAP (IN1 => n_13215, Y => a_N4186_aCLK);
dff_11706: DFF_a8237

    PORT MAP ( D => a_N4187_aD, CLK => a_N4187_aCLK, CLRN => vcc, PRN => vcc,
          Q => a_N4187);
xor2_11707: a_N4187_aD <=  n_13223  XOR n_13226;
or1_11708: n_13223 <=  n_13224;
and1_11709: n_13224 <=  n_13225;
delay_11710: n_13225  <= TRANSPORT a_N4186  ;
and1_11711: n_13226 <=  gnd;
delay_11712: n_13227  <= TRANSPORT clk  ;
filter_11713: FILTER_a8237

    PORT MAP (IN1 => n_13227, Y => a_N4187_aCLK);
delay_11714: a_N4170_aNOT  <= TRANSPORT a_EQ853  ;
xor2_11715: a_EQ853 <=  n_13231  XOR n_13236;
or2_11716: n_13231 <=  n_13232  OR n_13234;
and1_11717: n_13232 <=  n_13233;
delay_11718: n_13233  <= TRANSPORT a_N4187  ;
and1_11719: n_13234 <=  n_13235;
inv_11720: n_13235  <= TRANSPORT NOT a_N4186  ;
and1_11721: n_13236 <=  gnd;
dff_11722: DFF_a8237

    PORT MAP ( D => a_EQ866, CLK => a_SCHANNEL_F1_G_aCLK, CLRN => a_SCHANNEL_F1_G_aCLRN,
          PRN => vcc, Q => a_SCHANNEL_F1_G);
inv_11723: a_SCHANNEL_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11724: a_EQ866 <=  n_13243  XOR n_13252;
or2_11725: n_13243 <=  n_13244  OR n_13248;
and3_11726: n_13244 <=  n_13245  AND n_13246  AND n_13247;
delay_11727: n_13245  <= TRANSPORT a_N2563_aNOT  ;
delay_11728: n_13246  <= TRANSPORT a_LC4_B2  ;
inv_11729: n_13247  <= TRANSPORT NOT a_N4170_aNOT  ;
and3_11730: n_13248 <=  n_13249  AND n_13250  AND n_13251;
delay_11731: n_13249  <= TRANSPORT a_N2563_aNOT  ;
delay_11732: n_13250  <= TRANSPORT a_N4170_aNOT  ;
delay_11733: n_13251  <= TRANSPORT a_SCHANNEL_F1_G  ;
and1_11734: n_13252 <=  gnd;
delay_11735: n_13253  <= TRANSPORT clk  ;
filter_11736: FILTER_a8237

    PORT MAP (IN1 => n_13253, Y => a_SCHANNEL_F1_G_aCLK);
delay_11737: a_LC8_B26  <= TRANSPORT a_EQ547  ;
xor2_11738: a_EQ547 <=  n_13257  XOR n_13266;
or4_11739: n_13257 <=  n_13258  OR n_13260  OR n_13262  OR n_13264;
and1_11740: n_13258 <=  n_13259;
inv_11741: n_13259  <= TRANSPORT NOT a_SCOMMANDREG_F4_G  ;
and1_11742: n_13260 <=  n_13261;
inv_11743: n_13261  <= TRANSPORT NOT a_N2377  ;
and1_11744: n_13262 <=  n_13263;
delay_11745: n_13263  <= TRANSPORT a_N59  ;
and1_11746: n_13264 <=  n_13265;
inv_11747: n_13265  <= TRANSPORT NOT a_N2376  ;
and1_11748: n_13266 <=  gnd;
delay_11749: a_LC7_B26_aNOT  <= TRANSPORT a_LC7_B26_aNOT_aIN  ;
xor2_11750: a_LC7_B26_aNOT_aIN <=  n_13269  XOR n_13273;
or1_11751: n_13269 <=  n_13270;
and2_11752: n_13270 <=  n_13271  AND n_13272;
delay_11753: n_13271  <= TRANSPORT a_N2376  ;
delay_11754: n_13272  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
and1_11755: n_13273 <=  gnd;
delay_11756: a_LC6_B26  <= TRANSPORT a_EQ549  ;
xor2_11757: a_EQ549 <=  n_13276  XOR n_13283;
or2_11758: n_13276 <=  n_13277  OR n_13280;
and2_11759: n_13277 <=  n_13278  AND n_13279;
delay_11760: n_13278  <= TRANSPORT a_N55  ;
delay_11761: n_13279  <= TRANSPORT a_LC8_B26  ;
and2_11762: n_13280 <=  n_13281  AND n_13282;
inv_11763: n_13281  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_11764: n_13282  <= TRANSPORT a_LC7_B26_aNOT  ;
and1_11765: n_13283 <=  gnd;
delay_11766: a_LC4_B26  <= TRANSPORT a_EQ550  ;
xor2_11767: a_EQ550 <=  n_13286  XOR n_13295;
or3_11768: n_13286 <=  n_13287  OR n_13290  OR n_13293;
and2_11769: n_13287 <=  n_13288  AND n_13289;
inv_11770: n_13288  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_11771: n_13289  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
and2_11772: n_13290 <=  n_13291  AND n_13292;
inv_11773: n_13291  <= TRANSPORT NOT a_N88_aNOT  ;
delay_11774: n_13292  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
and1_11775: n_13293 <=  n_13294;
delay_11776: n_13294  <= TRANSPORT a_N55  ;
and1_11777: n_13295 <=  gnd;
delay_11778: a_LC3_B26  <= TRANSPORT a_EQ551  ;
xor2_11779: a_EQ551 <=  n_13298  XOR n_13305;
or2_11780: n_13298 <=  n_13299  OR n_13302;
and2_11781: n_13299 <=  n_13300  AND n_13301;
delay_11782: n_13300  <= TRANSPORT a_N59  ;
delay_11783: n_13301  <= TRANSPORT a_LC4_B26  ;
and2_11784: n_13302 <=  n_13303  AND n_13304;
inv_11785: n_13303  <= TRANSPORT NOT a_N2376  ;
delay_11786: n_13304  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
and1_11787: n_13305 <=  gnd;
delay_11788: a_LC2_B26  <= TRANSPORT a_EQ552  ;
xor2_11789: a_EQ552 <=  n_13308  XOR n_13315;
or2_11790: n_13308 <=  n_13309  OR n_13312;
and2_11791: n_13309 <=  n_13310  AND n_13311;
delay_11792: n_13310  <= TRANSPORT a_N2536  ;
delay_11793: n_13311  <= TRANSPORT a_LC6_B26  ;
and2_11794: n_13312 <=  n_13313  AND n_13314;
delay_11795: n_13313  <= TRANSPORT a_N2534  ;
delay_11796: n_13314  <= TRANSPORT a_LC3_B26  ;
and1_11797: n_13315 <=  gnd;
dff_11798: DFF_a8237

    PORT MAP ( D => a_EQ865, CLK => a_SCHANNEL_F0_G_aCLK, CLRN => a_SCHANNEL_F0_G_aCLRN,
          PRN => vcc, Q => a_SCHANNEL_F0_G);
inv_11799: a_SCHANNEL_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11800: a_EQ865 <=  n_13322  XOR n_13331;
or2_11801: n_13322 <=  n_13323  OR n_13327;
and3_11802: n_13323 <=  n_13324  AND n_13325  AND n_13326;
delay_11803: n_13324  <= TRANSPORT a_N2563_aNOT  ;
inv_11804: n_13325  <= TRANSPORT NOT a_N4170_aNOT  ;
delay_11805: n_13326  <= TRANSPORT a_LC2_B26  ;
and3_11806: n_13327 <=  n_13328  AND n_13329  AND n_13330;
delay_11807: n_13328  <= TRANSPORT a_N2563_aNOT  ;
delay_11808: n_13329  <= TRANSPORT a_N4170_aNOT  ;
delay_11809: n_13330  <= TRANSPORT a_SCHANNEL_F0_G  ;
and1_11810: n_13331 <=  gnd;
delay_11811: n_13332  <= TRANSPORT clk  ;
filter_11812: FILTER_a8237

    PORT MAP (IN1 => n_13332, Y => a_SCHANNEL_F0_G_aCLK);
dff_11813: DFF_a8237

    PORT MAP ( D => startdma_aD, CLK => startdma_aCLK, CLRN => vcc, PRN => vcc,
          Q => startdma);
xor2_11814: startdma_aD <=  n_13339  XOR n_13342;
or1_11815: n_13339 <=  n_13340;
and1_11816: n_13340 <=  n_13341;
inv_11817: n_13341  <= TRANSPORT NOT a_N4170_aNOT  ;
and1_11818: n_13342 <=  gnd;
delay_11819: n_13343  <= TRANSPORT clk  ;
filter_11820: FILTER_a8237

    PORT MAP (IN1 => n_13343, Y => startdma_aCLK);
dff_11821: DFF_a8237

    PORT MAP ( D => a_EQ1128, CLK => a_SCOMMANDREG_F5_G_aCLK, CLRN => a_SCOMMANDREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SCOMMANDREG_F5_G);
inv_11822: a_SCOMMANDREG_F5_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11823: a_EQ1128 <=  n_13352  XOR n_13361;
or2_11824: n_13352 <=  n_13353  OR n_13357;
and3_11825: n_13353 <=  n_13354  AND n_13355  AND n_13356;
delay_11826: n_13354  <= TRANSPORT a_N2563_aNOT  ;
delay_11827: n_13355  <= TRANSPORT a_N2571_aNOT  ;
delay_11828: n_13356  <= TRANSPORT a_SCOMMANDREG_F5_G  ;
and3_11829: n_13357 <=  n_13358  AND n_13359  AND n_13360;
delay_11830: n_13358  <= TRANSPORT a_N2563_aNOT  ;
inv_11831: n_13359  <= TRANSPORT NOT a_N2571_aNOT  ;
delay_11832: n_13360  <= TRANSPORT dbin(5)  ;
and1_11833: n_13361 <=  gnd;
delay_11834: n_13362  <= TRANSPORT clk  ;
filter_11835: FILTER_a8237

    PORT MAP (IN1 => n_13362, Y => a_SCOMMANDREG_F5_G_aCLK);
delay_11836: a_LC6_B3  <= TRANSPORT a_EQ529  ;
xor2_11837: a_EQ529 <=  n_13366  XOR n_13374;
or2_11838: n_13366 <=  n_13367  OR n_13371;
and3_11839: n_13367 <=  n_13368  AND n_13369  AND n_13370;
inv_11840: n_13368  <= TRANSPORT NOT a_N2356  ;
inv_11841: n_13369  <= TRANSPORT NOT a_N2369_aNOT  ;
inv_11842: n_13370  <= TRANSPORT NOT ready  ;
and2_11843: n_13371 <=  n_13372  AND n_13373;
inv_11844: n_13372  <= TRANSPORT NOT a_N67_aNOT  ;
inv_11845: n_13373  <= TRANSPORT NOT ready  ;
and1_11846: n_13374 <=  gnd;
delay_11847: a_LC7_B16  <= TRANSPORT a_LC7_B16_aIN  ;
xor2_11848: a_LC7_B16_aIN <=  n_13377  XOR n_13382;
or1_11849: n_13377 <=  n_13378;
and3_11850: n_13378 <=  n_13379  AND n_13380  AND n_13381;
delay_11851: n_13379  <= TRANSPORT a_N820  ;
inv_11852: n_13380  <= TRANSPORT NOT a_N822  ;
inv_11853: n_13381  <= TRANSPORT NOT a_N823  ;
and1_11854: n_13382 <=  gnd;
delay_11855: a_LC8_B16  <= TRANSPORT a_EQ531  ;
xor2_11856: a_EQ531 <=  n_13385  XOR n_13394;
or3_11857: n_13385 <=  n_13386  OR n_13389  OR n_13392;
and2_11858: n_13386 <=  n_13387  AND n_13388;
delay_11859: n_13387  <= TRANSPORT a_N2359_aNOT  ;
inv_11860: n_13388  <= TRANSPORT NOT startdma  ;
and2_11861: n_13389 <=  n_13390  AND n_13391;
delay_11862: n_13390  <= TRANSPORT a_N2591  ;
delay_11863: n_13391  <= TRANSPORT a_N2359_aNOT  ;
and1_11864: n_13392 <=  n_13393;
delay_11865: n_13393  <= TRANSPORT a_LC7_B16  ;
and1_11866: n_13394 <=  gnd;
delay_11867: a_LC1_B2  <= TRANSPORT a_LC1_B2_aIN  ;
xor2_11868: a_LC1_B2_aIN <=  n_13397  XOR n_13402;
or1_11869: n_13397 <=  n_13398;
and3_11870: n_13398 <=  n_13399  AND n_13400  AND n_13401;
inv_11871: n_13399  <= TRANSPORT NOT a_N1566  ;
inv_11872: n_13400  <= TRANSPORT NOT a_SCOMMANDREG_F2_G  ;
inv_11873: n_13401  <= TRANSPORT NOT a_N823  ;
and1_11874: n_13402 <=  gnd;
delay_11875: a_N1381  <= TRANSPORT a_EQ428  ;
xor2_11876: a_EQ428 <=  n_13405  XOR n_13415;
or3_11877: n_13405 <=  n_13406  OR n_13409  OR n_13412;
and2_11878: n_13406 <=  n_13407  AND n_13408;
delay_11879: n_13407  <= TRANSPORT a_N2536  ;
delay_11880: n_13408  <= TRANSPORT a_LC1_B2  ;
and2_11881: n_13409 <=  n_13410  AND n_13411;
inv_11882: n_13410  <= TRANSPORT NOT a_N55  ;
delay_11883: n_13411  <= TRANSPORT a_LC1_B2  ;
and2_11884: n_13412 <=  n_13413  AND n_13414;
delay_11885: n_13413  <= TRANSPORT a_N2606  ;
delay_11886: n_13414  <= TRANSPORT a_LC1_B2  ;
and1_11887: n_13415 <=  gnd;
delay_11888: a_LC7_B3  <= TRANSPORT a_EQ532  ;
xor2_11889: a_EQ532 <=  n_13418  XOR n_13427;
or4_11890: n_13418 <=  n_13419  OR n_13421  OR n_13423  OR n_13425;
and1_11891: n_13419 <=  n_13420;
delay_11892: n_13420  <= TRANSPORT a_LC6_B3  ;
and1_11893: n_13421 <=  n_13422;
delay_11894: n_13422  <= TRANSPORT a_LC8_B16  ;
and1_11895: n_13423 <=  n_13424;
delay_11896: n_13424  <= TRANSPORT a_N1381  ;
and1_11897: n_13425 <=  n_13426;
delay_11898: n_13426  <= TRANSPORT a_LC4_B13  ;
and1_11899: n_13427 <=  gnd;
delay_11900: a_LC2_F17  <= TRANSPORT a_EQ526  ;
xor2_11901: a_EQ526 <=  n_13430  XOR n_13439;
or4_11902: n_13430 <=  n_13431  OR n_13433  OR n_13435  OR n_13437;
and1_11903: n_13431 <=  n_13432;
inv_11904: n_13432  <= TRANSPORT NOT a_LC1_C16  ;
and1_11905: n_13433 <=  n_13434;
inv_11906: n_13434  <= TRANSPORT NOT a_LC5_D27  ;
and1_11907: n_13435 <=  n_13436;
inv_11908: n_13436  <= TRANSPORT NOT a_LC3_F6  ;
and1_11909: n_13437 <=  n_13438;
inv_11910: n_13438  <= TRANSPORT NOT a_LC2_C24  ;
and1_11911: n_13439 <=  gnd;
delay_11912: a_LC1_F17  <= TRANSPORT a_EQ527  ;
xor2_11913: a_EQ527 <=  n_13442  XOR n_13451;
or4_11914: n_13442 <=  n_13443  OR n_13445  OR n_13447  OR n_13449;
and1_11915: n_13443 <=  n_13444;
inv_11916: n_13444  <= TRANSPORT NOT a_LC4_C16  ;
and1_11917: n_13445 <=  n_13446;
inv_11918: n_13446  <= TRANSPORT NOT a_LC7_C17  ;
and1_11919: n_13447 <=  n_13448;
inv_11920: n_13448  <= TRANSPORT NOT a_LC7_D18  ;
and1_11921: n_13449 <=  n_13450;
delay_11922: n_13450  <= TRANSPORT a_LC2_F17  ;
and1_11923: n_13451 <=  gnd;
delay_11924: a_LC6_F17  <= TRANSPORT a_EQ524  ;
xor2_11925: a_EQ524 <=  n_13454  XOR n_13463;
or4_11926: n_13454 <=  n_13455  OR n_13457  OR n_13459  OR n_13461;
and1_11927: n_13455 <=  n_13456;
delay_11928: n_13456  <= TRANSPORT a_LC1_C16  ;
and1_11929: n_13457 <=  n_13458;
delay_11930: n_13458  <= TRANSPORT a_LC7_C17  ;
and1_11931: n_13459 <=  n_13460;
delay_11932: n_13460  <= TRANSPORT a_LC5_D27  ;
and1_11933: n_13461 <=  n_13462;
delay_11934: n_13462  <= TRANSPORT a_LC2_C24  ;
and1_11935: n_13463 <=  gnd;
delay_11936: a_LC4_F17  <= TRANSPORT a_EQ525  ;
xor2_11937: a_EQ525 <=  n_13466  XOR n_13475;
or4_11938: n_13466 <=  n_13467  OR n_13469  OR n_13471  OR n_13473;
and1_11939: n_13467 <=  n_13468;
delay_11940: n_13468  <= TRANSPORT a_LC6_F17  ;
and1_11941: n_13469 <=  n_13470;
delay_11942: n_13470  <= TRANSPORT a_LC7_D18  ;
and1_11943: n_13471 <=  n_13472;
delay_11944: n_13472  <= TRANSPORT a_LC3_F6  ;
and1_11945: n_13473 <=  n_13474;
delay_11946: n_13474  <= TRANSPORT a_LC4_C16  ;
and1_11947: n_13475 <=  gnd;
delay_11948: a_LC5_F17  <= TRANSPORT a_EQ528  ;
xor2_11949: a_EQ528 <=  n_13478  XOR n_13491;
or4_11950: n_13478 <=  n_13479  OR n_13482  OR n_13485  OR n_13488;
and2_11951: n_13479 <=  n_13480  AND n_13481;
delay_11952: n_13480  <= TRANSPORT a_LC1_F17  ;
delay_11953: n_13481  <= TRANSPORT a_LC4_F10  ;
and2_11954: n_13482 <=  n_13483  AND n_13484;
inv_11955: n_13483  <= TRANSPORT NOT a_N2529  ;
delay_11956: n_13484  <= TRANSPORT a_LC4_F10  ;
and2_11957: n_13485 <=  n_13486  AND n_13487;
delay_11958: n_13486  <= TRANSPORT a_LC4_F17  ;
inv_11959: n_13487  <= TRANSPORT NOT a_LC4_F10  ;
and2_11960: n_13488 <=  n_13489  AND n_13490;
delay_11961: n_13489  <= TRANSPORT a_N2529  ;
inv_11962: n_13490  <= TRANSPORT NOT a_LC4_F10  ;
and1_11963: n_13491 <=  gnd;
dff_11964: DFF_a8237

    PORT MAP ( D => a_EQ309, CLK => a_N823_aCLK, CLRN => a_N823_aCLRN, PRN => vcc,
          Q => a_N823);
inv_11965: a_N823_aCLRN  <= TRANSPORT NOT reset  ;
xor2_11966: a_EQ309 <=  n_13498  XOR n_13506;
or2_11967: n_13498 <=  n_13499  OR n_13502;
and2_11968: n_13499 <=  n_13500  AND n_13501;
delay_11969: n_13500  <= TRANSPORT a_N2563_aNOT  ;
delay_11970: n_13501  <= TRANSPORT a_LC7_B3  ;
and3_11971: n_13502 <=  n_13503  AND n_13504  AND n_13505;
delay_11972: n_13503  <= TRANSPORT a_N2563_aNOT  ;
delay_11973: n_13504  <= TRANSPORT a_N2394  ;
delay_11974: n_13505  <= TRANSPORT a_LC5_F17  ;
and1_11975: n_13506 <=  gnd;
delay_11976: n_13507  <= TRANSPORT clk  ;
filter_11977: FILTER_a8237

    PORT MAP (IN1 => n_13507, Y => a_N823_aCLK);
delay_11978: a_LC1_D18  <= TRANSPORT a_EQ450  ;
xor2_11979: a_EQ450 <=  n_13511  XOR n_13518;
or2_11980: n_13511 <=  n_13512  OR n_13515;
and2_11981: n_13512 <=  n_13513  AND n_13514;
inv_11982: n_13513  <= TRANSPORT NOT a_N2376  ;
delay_11983: n_13514  <= TRANSPORT a_SCH2ADDRREG_F0_G  ;
and2_11984: n_13515 <=  n_13516  AND n_13517;
inv_11985: n_13516  <= TRANSPORT NOT a_N2377  ;
delay_11986: n_13517  <= TRANSPORT a_SCH3ADDRREG_F0_G  ;
and1_11987: n_13518 <=  gnd;
delay_11988: a_LC4_D18  <= TRANSPORT a_EQ453  ;
xor2_11989: a_EQ453 <=  n_13521  XOR n_13537;
or4_11990: n_13521 <=  n_13522  OR n_13526  OR n_13530  OR n_13534;
and3_11991: n_13522 <=  n_13523  AND n_13524  AND n_13525;
delay_11992: n_13523  <= TRANSPORT a_N2557  ;
inv_11993: n_13524  <= TRANSPORT NOT a_SCOMMANDREG_F1_G  ;
inv_11994: n_13525  <= TRANSPORT NOT a_LC7_D18  ;
and3_11995: n_13526 <=  n_13527  AND n_13528  AND n_13529;
delay_11996: n_13527  <= TRANSPORT a_N2557  ;
delay_11997: n_13528  <= TRANSPORT a_N2598_aNOT  ;
inv_11998: n_13529  <= TRANSPORT NOT a_LC7_D18  ;
and3_11999: n_13530 <=  n_13531  AND n_13532  AND n_13533;
inv_12000: n_13531  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12001: n_13532  <= TRANSPORT a_SCOMMANDREG_F1_G  ;
delay_12002: n_13533  <= TRANSPORT a_LC7_D18  ;
and2_12003: n_13534 <=  n_13535  AND n_13536;
inv_12004: n_13535  <= TRANSPORT NOT a_N2557  ;
delay_12005: n_13536  <= TRANSPORT a_LC7_D18  ;
and1_12006: n_13537 <=  gnd;
delay_12007: a_N1486  <= TRANSPORT a_EQ454  ;
xor2_12008: a_EQ454 <=  n_13540  XOR n_13547;
or2_12009: n_13540 <=  n_13541  OR n_13544;
and2_12010: n_13541 <=  n_13542  AND n_13543;
delay_12011: n_13542  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12012: n_13543  <= TRANSPORT a_SCH1ADDRREG_F0_G  ;
and2_12013: n_13544 <=  n_13545  AND n_13546;
inv_12014: n_13545  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12015: n_13546  <= TRANSPORT a_SCH0ADDRREG_F0_G  ;
and1_12016: n_13547 <=  gnd;
delay_12017: a_N1471  <= TRANSPORT a_EQ452  ;
xor2_12018: a_EQ452 <=  n_13550  XOR n_13559;
or3_12019: n_13550 <=  n_13551  OR n_13554  OR n_13557;
and2_12020: n_13551 <=  n_13552  AND n_13553;
inv_12021: n_13552  <= TRANSPORT NOT a_N2531  ;
delay_12022: n_13553  <= TRANSPORT a_LC4_D18  ;
and2_12023: n_13554 <=  n_13555  AND n_13556;
delay_12024: n_13555  <= TRANSPORT a_N2531  ;
delay_12025: n_13556  <= TRANSPORT a_N1486  ;
and1_12026: n_13557 <=  n_13558;
delay_12027: n_13558  <= TRANSPORT startdma  ;
and1_12028: n_13559 <=  gnd;
delay_12029: a_LC2_D18  <= TRANSPORT a_EQ451  ;
xor2_12030: a_EQ451 <=  n_13562  XOR n_13569;
or2_12031: n_13562 <=  n_13563  OR n_13566;
and2_12032: n_13563 <=  n_13564  AND n_13565;
inv_12033: n_13564  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12034: n_13565  <= TRANSPORT a_SCH0ADDRREG_F0_G  ;
and2_12035: n_13566 <=  n_13567  AND n_13568;
inv_12036: n_13567  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12037: n_13568  <= TRANSPORT a_SCH1ADDRREG_F0_G  ;
and1_12038: n_13569 <=  gnd;
dff_12039: DFF_a8237

    PORT MAP ( D => a_EQ044, CLK => a_LC7_D18_aCLK, CLRN => a_LC7_D18_aCLRN,
          PRN => vcc, Q => a_LC7_D18);
inv_12040: a_LC7_D18_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12041: a_EQ044 <=  n_13576  XOR n_13586;
or3_12042: n_13576 <=  n_13577  OR n_13580  OR n_13583;
and2_12043: n_13577 <=  n_13578  AND n_13579;
delay_12044: n_13578  <= TRANSPORT a_LC1_D18  ;
delay_12045: n_13579  <= TRANSPORT a_N1471  ;
and2_12046: n_13580 <=  n_13581  AND n_13582;
delay_12047: n_13581  <= TRANSPORT a_N1471  ;
delay_12048: n_13582  <= TRANSPORT a_LC2_D18  ;
and2_12049: n_13583 <=  n_13584  AND n_13585;
inv_12050: n_13584  <= TRANSPORT NOT startdma  ;
delay_12051: n_13585  <= TRANSPORT a_N1471  ;
and1_12052: n_13586 <=  gnd;
delay_12053: n_13587  <= TRANSPORT clk  ;
filter_12054: FILTER_a8237

    PORT MAP (IN1 => n_13587, Y => a_LC7_D18_aCLK);
delay_12055: a_LC4_C17  <= TRANSPORT a_EQ523  ;
xor2_12056: a_EQ523 <=  n_13591  XOR n_13602;
or3_12057: n_13591 <=  n_13592  OR n_13596  OR n_13599;
and3_12058: n_13592 <=  n_13593  AND n_13594  AND n_13595;
delay_12059: n_13593  <= TRANSPORT a_N2557  ;
delay_12060: n_13594  <= TRANSPORT a_N2530_aNOT  ;
delay_12061: n_13595  <= TRANSPORT a_N3059  ;
and2_12062: n_13596 <=  n_13597  AND n_13598;
inv_12063: n_13597  <= TRANSPORT NOT a_N2530_aNOT  ;
delay_12064: n_13598  <= TRANSPORT a_LC7_C17  ;
and2_12065: n_13599 <=  n_13600  AND n_13601;
inv_12066: n_13600  <= TRANSPORT NOT a_N2557  ;
delay_12067: n_13601  <= TRANSPORT a_LC7_C17  ;
and1_12068: n_13602 <=  gnd;
delay_12069: a_N1904  <= TRANSPORT a_EQ519  ;
xor2_12070: a_EQ519 <=  n_13605  XOR n_13612;
or2_12071: n_13605 <=  n_13606  OR n_13609;
and2_12072: n_13606 <=  n_13607  AND n_13608;
delay_12073: n_13607  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12074: n_13608  <= TRANSPORT a_SCH1ADDRREG_F1_G  ;
and2_12075: n_13609 <=  n_13610  AND n_13611;
inv_12076: n_13610  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12077: n_13611  <= TRANSPORT a_SCH0ADDRREG_F1_G  ;
and1_12078: n_13612 <=  gnd;
delay_12079: a_LC5_C17  <= TRANSPORT a_EQ522  ;
xor2_12080: a_EQ522 <=  n_13615  XOR n_13622;
or2_12081: n_13615 <=  n_13616  OR n_13619;
and2_12082: n_13616 <=  n_13617  AND n_13618;
inv_12083: n_13617  <= TRANSPORT NOT a_N2531  ;
delay_12084: n_13618  <= TRANSPORT a_LC4_C17  ;
and2_12085: n_13619 <=  n_13620  AND n_13621;
delay_12086: n_13620  <= TRANSPORT a_N2531  ;
delay_12087: n_13621  <= TRANSPORT a_N1904  ;
and1_12088: n_13622 <=  gnd;
delay_12089: a_LC2_C17  <= TRANSPORT a_EQ521  ;
xor2_12090: a_EQ521 <=  n_13625  XOR n_13632;
or2_12091: n_13625 <=  n_13626  OR n_13629;
and2_12092: n_13626 <=  n_13627  AND n_13628;
inv_12093: n_13627  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12094: n_13628  <= TRANSPORT a_SCH1ADDRREG_F1_G  ;
and2_12095: n_13629 <=  n_13630  AND n_13631;
inv_12096: n_13630  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12097: n_13631  <= TRANSPORT a_SCH0ADDRREG_F1_G  ;
and1_12098: n_13632 <=  gnd;
delay_12099: a_LC1_C17  <= TRANSPORT a_EQ520  ;
xor2_12100: a_EQ520 <=  n_13635  XOR n_13642;
or2_12101: n_13635 <=  n_13636  OR n_13639;
and2_12102: n_13636 <=  n_13637  AND n_13638;
inv_12103: n_13637  <= TRANSPORT NOT a_N2376  ;
delay_12104: n_13638  <= TRANSPORT a_SCH2ADDRREG_F1_G  ;
and2_12105: n_13639 <=  n_13640  AND n_13641;
inv_12106: n_13640  <= TRANSPORT NOT a_N2377  ;
delay_12107: n_13641  <= TRANSPORT a_SCH3ADDRREG_F1_G  ;
and1_12108: n_13642 <=  gnd;
dff_12109: DFF_a8237

    PORT MAP ( D => a_EQ043, CLK => a_LC7_C17_aCLK, CLRN => a_LC7_C17_aCLRN,
          PRN => vcc, Q => a_LC7_C17);
inv_12110: a_LC7_C17_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12111: a_EQ043 <=  n_13649  XOR n_13659;
or3_12112: n_13649 <=  n_13650  OR n_13653  OR n_13656;
and2_12113: n_13650 <=  n_13651  AND n_13652;
inv_12114: n_13651  <= TRANSPORT NOT startdma  ;
delay_12115: n_13652  <= TRANSPORT a_LC5_C17  ;
and2_12116: n_13653 <=  n_13654  AND n_13655;
delay_12117: n_13654  <= TRANSPORT startdma  ;
delay_12118: n_13655  <= TRANSPORT a_LC2_C17  ;
and2_12119: n_13656 <=  n_13657  AND n_13658;
delay_12120: n_13657  <= TRANSPORT startdma  ;
delay_12121: n_13658  <= TRANSPORT a_LC1_C17  ;
and1_12122: n_13659 <=  gnd;
delay_12123: n_13660  <= TRANSPORT clk  ;
filter_12124: FILTER_a8237

    PORT MAP (IN1 => n_13660, Y => a_LC7_C17_aCLK);
delay_12125: a_N1337_aNOT  <= TRANSPORT a_EQ424  ;
xor2_12126: a_EQ424 <=  n_13664  XOR n_13671;
or2_12127: n_13664 <=  n_13665  OR n_13668;
and2_12128: n_13665 <=  n_13666  AND n_13667;
delay_12129: n_13666  <= TRANSPORT a_N2557  ;
delay_12130: n_13667  <= TRANSPORT a_N2542  ;
and2_12131: n_13668 <=  n_13669  AND n_13670;
inv_12132: n_13669  <= TRANSPORT NOT a_N2557  ;
delay_12133: n_13670  <= TRANSPORT a_LC4_C16  ;
and1_12134: n_13671 <=  gnd;
delay_12135: a_N1321  <= TRANSPORT a_EQ413  ;
xor2_12136: a_EQ413 <=  n_13674  XOR n_13681;
or2_12137: n_13674 <=  n_13675  OR n_13678;
and2_12138: n_13675 <=  n_13676  AND n_13677;
delay_12139: n_13676  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12140: n_13677  <= TRANSPORT a_SCH1ADDRREG_F2_G  ;
and2_12141: n_13678 <=  n_13679  AND n_13680;
inv_12142: n_13679  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12143: n_13680  <= TRANSPORT a_SCH0ADDRREG_F2_G  ;
and1_12144: n_13681 <=  gnd;
delay_12145: a_LC8_C16  <= TRANSPORT a_EQ412  ;
xor2_12146: a_EQ412 <=  n_13684  XOR n_13691;
or2_12147: n_13684 <=  n_13685  OR n_13688;
and2_12148: n_13685 <=  n_13686  AND n_13687;
inv_12149: n_13686  <= TRANSPORT NOT a_N2531  ;
delay_12150: n_13687  <= TRANSPORT a_N1337_aNOT  ;
and2_12151: n_13688 <=  n_13689  AND n_13690;
delay_12152: n_13689  <= TRANSPORT a_N2531  ;
delay_12153: n_13690  <= TRANSPORT a_N1321  ;
and1_12154: n_13691 <=  gnd;
delay_12155: a_LC2_C16  <= TRANSPORT a_EQ415  ;
xor2_12156: a_EQ415 <=  n_13694  XOR n_13701;
or2_12157: n_13694 <=  n_13695  OR n_13698;
and2_12158: n_13695 <=  n_13696  AND n_13697;
inv_12159: n_13696  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12160: n_13697  <= TRANSPORT a_SCH1ADDRREG_F2_G  ;
and2_12161: n_13698 <=  n_13699  AND n_13700;
inv_12162: n_13699  <= TRANSPORT NOT a_N2377  ;
delay_12163: n_13700  <= TRANSPORT a_SCH3ADDRREG_F2_G  ;
and1_12164: n_13701 <=  gnd;
delay_12165: a_LC5_C16  <= TRANSPORT a_EQ414  ;
xor2_12166: a_EQ414 <=  n_13704  XOR n_13711;
or2_12167: n_13704 <=  n_13705  OR n_13708;
and2_12168: n_13705 <=  n_13706  AND n_13707;
inv_12169: n_13706  <= TRANSPORT NOT a_N2376  ;
delay_12170: n_13707  <= TRANSPORT a_SCH2ADDRREG_F2_G  ;
and2_12171: n_13708 <=  n_13709  AND n_13710;
inv_12172: n_13709  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12173: n_13710  <= TRANSPORT a_SCH0ADDRREG_F2_G  ;
and1_12174: n_13711 <=  gnd;
dff_12175: DFF_a8237

    PORT MAP ( D => a_EQ042, CLK => a_LC4_C16_aCLK, CLRN => a_LC4_C16_aCLRN,
          PRN => vcc, Q => a_LC4_C16);
inv_12176: a_LC4_C16_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12177: a_EQ042 <=  n_13718  XOR n_13728;
or3_12178: n_13718 <=  n_13719  OR n_13722  OR n_13725;
and2_12179: n_13719 <=  n_13720  AND n_13721;
inv_12180: n_13720  <= TRANSPORT NOT startdma  ;
delay_12181: n_13721  <= TRANSPORT a_LC8_C16  ;
and2_12182: n_13722 <=  n_13723  AND n_13724;
delay_12183: n_13723  <= TRANSPORT startdma  ;
delay_12184: n_13724  <= TRANSPORT a_LC2_C16  ;
and2_12185: n_13725 <=  n_13726  AND n_13727;
delay_12186: n_13726  <= TRANSPORT startdma  ;
delay_12187: n_13727  <= TRANSPORT a_LC5_C16  ;
and1_12188: n_13728 <=  gnd;
delay_12189: n_13729  <= TRANSPORT clk  ;
filter_12190: FILTER_a8237

    PORT MAP (IN1 => n_13729, Y => a_LC4_C16_aCLK);
delay_12191: a_LC5_C24  <= TRANSPORT a_EQ289  ;
xor2_12192: a_EQ289 <=  n_13733  XOR n_13740;
or2_12193: n_13733 <=  n_13734  OR n_13737;
and2_12194: n_13734 <=  n_13735  AND n_13736;
delay_12195: n_13735  <= TRANSPORT a_N2557  ;
delay_12196: n_13736  <= TRANSPORT a_N2543  ;
and2_12197: n_13737 <=  n_13738  AND n_13739;
inv_12198: n_13738  <= TRANSPORT NOT a_N2557  ;
delay_12199: n_13739  <= TRANSPORT a_LC2_C24  ;
and1_12200: n_13740 <=  gnd;
delay_12201: a_LC6_C24  <= TRANSPORT a_EQ290  ;
xor2_12202: a_EQ290 <=  n_13743  XOR n_13750;
or2_12203: n_13743 <=  n_13744  OR n_13747;
and2_12204: n_13744 <=  n_13745  AND n_13746;
delay_12205: n_13745  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12206: n_13746  <= TRANSPORT a_SCH1ADDRREG_F3_G  ;
and2_12207: n_13747 <=  n_13748  AND n_13749;
inv_12208: n_13748  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12209: n_13749  <= TRANSPORT a_SCH0ADDRREG_F3_G  ;
and1_12210: n_13750 <=  gnd;
delay_12211: a_N725_aNOT  <= TRANSPORT a_EQ291  ;
xor2_12212: a_EQ291 <=  n_13753  XOR n_13760;
or2_12213: n_13753 <=  n_13754  OR n_13757;
and2_12214: n_13754 <=  n_13755  AND n_13756;
inv_12215: n_13755  <= TRANSPORT NOT a_N2531  ;
delay_12216: n_13756  <= TRANSPORT a_LC5_C24  ;
and2_12217: n_13757 <=  n_13758  AND n_13759;
delay_12218: n_13758  <= TRANSPORT a_N2531  ;
delay_12219: n_13759  <= TRANSPORT a_LC6_C24  ;
and1_12220: n_13760 <=  gnd;
delay_12221: a_LC4_C24  <= TRANSPORT a_EQ293  ;
xor2_12222: a_EQ293 <=  n_13763  XOR n_13770;
or2_12223: n_13763 <=  n_13764  OR n_13767;
and2_12224: n_13764 <=  n_13765  AND n_13766;
inv_12225: n_13765  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12226: n_13766  <= TRANSPORT a_SCH0ADDRREG_F3_G  ;
and2_12227: n_13767 <=  n_13768  AND n_13769;
inv_12228: n_13768  <= TRANSPORT NOT a_N2376  ;
delay_12229: n_13769  <= TRANSPORT a_SCH2ADDRREG_F3_G  ;
and1_12230: n_13770 <=  gnd;
delay_12231: a_LC3_C24  <= TRANSPORT a_EQ292  ;
xor2_12232: a_EQ292 <=  n_13773  XOR n_13780;
or2_12233: n_13773 <=  n_13774  OR n_13777;
and2_12234: n_13774 <=  n_13775  AND n_13776;
inv_12235: n_13775  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12236: n_13776  <= TRANSPORT a_SCH1ADDRREG_F3_G  ;
and2_12237: n_13777 <=  n_13778  AND n_13779;
inv_12238: n_13778  <= TRANSPORT NOT a_N2377  ;
delay_12239: n_13779  <= TRANSPORT a_SCH3ADDRREG_F3_G  ;
and1_12240: n_13780 <=  gnd;
dff_12241: DFF_a8237

    PORT MAP ( D => a_EQ041, CLK => a_LC2_C24_aCLK, CLRN => a_LC2_C24_aCLRN,
          PRN => vcc, Q => a_LC2_C24);
inv_12242: a_LC2_C24_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12243: a_EQ041 <=  n_13787  XOR n_13797;
or3_12244: n_13787 <=  n_13788  OR n_13791  OR n_13794;
and2_12245: n_13788 <=  n_13789  AND n_13790;
inv_12246: n_13789  <= TRANSPORT NOT startdma  ;
delay_12247: n_13790  <= TRANSPORT a_N725_aNOT  ;
and2_12248: n_13791 <=  n_13792  AND n_13793;
delay_12249: n_13792  <= TRANSPORT startdma  ;
delay_12250: n_13793  <= TRANSPORT a_LC4_C24  ;
and2_12251: n_13794 <=  n_13795  AND n_13796;
delay_12252: n_13795  <= TRANSPORT startdma  ;
delay_12253: n_13796  <= TRANSPORT a_LC3_C24  ;
and1_12254: n_13797 <=  gnd;
delay_12255: n_13798  <= TRANSPORT clk  ;
filter_12256: FILTER_a8237

    PORT MAP (IN1 => n_13798, Y => a_LC2_C24_aCLK);
delay_12257: a_N1725_aNOT  <= TRANSPORT a_EQ495  ;
xor2_12258: a_EQ495 <=  n_13802  XOR n_13809;
or2_12259: n_13802 <=  n_13803  OR n_13806;
and2_12260: n_13803 <=  n_13804  AND n_13805;
delay_12261: n_13804  <= TRANSPORT a_N2557  ;
delay_12262: n_13805  <= TRANSPORT a_N2544  ;
and2_12263: n_13806 <=  n_13807  AND n_13808;
inv_12264: n_13807  <= TRANSPORT NOT a_N2557  ;
delay_12265: n_13808  <= TRANSPORT a_LC1_C16  ;
and1_12266: n_13809 <=  gnd;
delay_12267: a_N1729  <= TRANSPORT a_EQ497  ;
xor2_12268: a_EQ497 <=  n_13812  XOR n_13819;
or2_12269: n_13812 <=  n_13813  OR n_13816;
and2_12270: n_13813 <=  n_13814  AND n_13815;
inv_12271: n_13814  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12272: n_13815  <= TRANSPORT a_SCH0ADDRREG_F4_G  ;
and2_12273: n_13816 <=  n_13817  AND n_13818;
delay_12274: n_13817  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12275: n_13818  <= TRANSPORT a_SCH1ADDRREG_F4_G  ;
and1_12276: n_13819 <=  gnd;
delay_12277: a_LC3_C15  <= TRANSPORT a_EQ489  ;
xor2_12278: a_EQ489 <=  n_13822  XOR n_13829;
or2_12279: n_13822 <=  n_13823  OR n_13826;
and2_12280: n_13823 <=  n_13824  AND n_13825;
inv_12281: n_13824  <= TRANSPORT NOT a_N2531  ;
delay_12282: n_13825  <= TRANSPORT a_N1725_aNOT  ;
and2_12283: n_13826 <=  n_13827  AND n_13828;
delay_12284: n_13827  <= TRANSPORT a_N2531  ;
delay_12285: n_13828  <= TRANSPORT a_N1729  ;
and1_12286: n_13829 <=  gnd;
delay_12287: a_LC3_C16  <= TRANSPORT a_EQ491  ;
xor2_12288: a_EQ491 <=  n_13832  XOR n_13839;
or2_12289: n_13832 <=  n_13833  OR n_13836;
and2_12290: n_13833 <=  n_13834  AND n_13835;
inv_12291: n_13834  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12292: n_13835  <= TRANSPORT a_SCH1ADDRREG_F4_G  ;
and2_12293: n_13836 <=  n_13837  AND n_13838;
inv_12294: n_13837  <= TRANSPORT NOT a_N2376  ;
delay_12295: n_13838  <= TRANSPORT a_SCH2ADDRREG_F4_G  ;
and1_12296: n_13839 <=  gnd;
delay_12297: a_LC4_C22  <= TRANSPORT a_EQ490  ;
xor2_12298: a_EQ490 <=  n_13842  XOR n_13849;
or2_12299: n_13842 <=  n_13843  OR n_13846;
and2_12300: n_13843 <=  n_13844  AND n_13845;
inv_12301: n_13844  <= TRANSPORT NOT a_N2377  ;
delay_12302: n_13845  <= TRANSPORT a_SCH3ADDRREG_F4_G  ;
and2_12303: n_13846 <=  n_13847  AND n_13848;
inv_12304: n_13847  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12305: n_13848  <= TRANSPORT a_SCH0ADDRREG_F4_G  ;
and1_12306: n_13849 <=  gnd;
dff_12307: DFF_a8237

    PORT MAP ( D => a_EQ040, CLK => a_LC1_C16_aCLK, CLRN => a_LC1_C16_aCLRN,
          PRN => vcc, Q => a_LC1_C16);
inv_12308: a_LC1_C16_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12309: a_EQ040 <=  n_13856  XOR n_13866;
or3_12310: n_13856 <=  n_13857  OR n_13860  OR n_13863;
and2_12311: n_13857 <=  n_13858  AND n_13859;
inv_12312: n_13858  <= TRANSPORT NOT startdma  ;
delay_12313: n_13859  <= TRANSPORT a_LC3_C15  ;
and2_12314: n_13860 <=  n_13861  AND n_13862;
delay_12315: n_13861  <= TRANSPORT startdma  ;
delay_12316: n_13862  <= TRANSPORT a_LC3_C16  ;
and2_12317: n_13863 <=  n_13864  AND n_13865;
delay_12318: n_13864  <= TRANSPORT startdma  ;
delay_12319: n_13865  <= TRANSPORT a_LC4_C22  ;
and1_12320: n_13866 <=  gnd;
delay_12321: n_13867  <= TRANSPORT clk  ;
filter_12322: FILTER_a8237

    PORT MAP (IN1 => n_13867, Y => a_LC1_C16_aCLK);
delay_12323: a_LC6_F6  <= TRANSPORT a_EQ237  ;
xor2_12324: a_EQ237 <=  n_13871  XOR n_13878;
or2_12325: n_13871 <=  n_13872  OR n_13875;
and2_12326: n_13872 <=  n_13873  AND n_13874;
delay_12327: n_13873  <= TRANSPORT a_N2557  ;
delay_12328: n_13874  <= TRANSPORT a_N2545  ;
and2_12329: n_13875 <=  n_13876  AND n_13877;
inv_12330: n_13876  <= TRANSPORT NOT a_N2557  ;
delay_12331: n_13877  <= TRANSPORT a_LC3_F6  ;
and1_12332: n_13878 <=  gnd;
delay_12333: a_LC5_F6  <= TRANSPORT a_EQ238  ;
xor2_12334: a_EQ238 <=  n_13881  XOR n_13888;
or2_12335: n_13881 <=  n_13882  OR n_13885;
and2_12336: n_13882 <=  n_13883  AND n_13884;
inv_12337: n_13883  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12338: n_13884  <= TRANSPORT a_SCH0ADDRREG_F5_G  ;
and2_12339: n_13885 <=  n_13886  AND n_13887;
delay_12340: n_13886  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12341: n_13887  <= TRANSPORT a_SCH1ADDRREG_F5_G  ;
and1_12342: n_13888 <=  gnd;
delay_12343: a_N423_aNOT  <= TRANSPORT a_EQ241  ;
xor2_12344: a_EQ241 <=  n_13891  XOR n_13902;
or3_12345: n_13891 <=  n_13892  OR n_13895  OR n_13898;
and2_12346: n_13892 <=  n_13893  AND n_13894;
inv_12347: n_13893  <= TRANSPORT NOT a_N2557  ;
delay_12348: n_13894  <= TRANSPORT a_LC6_F6  ;
and2_12349: n_13895 <=  n_13896  AND n_13897;
inv_12350: n_13896  <= TRANSPORT NOT a_N2591  ;
delay_12351: n_13897  <= TRANSPORT a_LC6_F6  ;
and3_12352: n_13898 <=  n_13899  AND n_13900  AND n_13901;
delay_12353: n_13899  <= TRANSPORT a_N2557  ;
delay_12354: n_13900  <= TRANSPORT a_N2591  ;
delay_12355: n_13901  <= TRANSPORT a_LC5_F6  ;
and1_12356: n_13902 <=  gnd;
delay_12357: a_LC2_F6  <= TRANSPORT a_EQ240  ;
xor2_12358: a_EQ240 <=  n_13905  XOR n_13912;
or2_12359: n_13905 <=  n_13906  OR n_13909;
and2_12360: n_13906 <=  n_13907  AND n_13908;
inv_12361: n_13907  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12362: n_13908  <= TRANSPORT a_SCH1ADDRREG_F5_G  ;
and2_12363: n_13909 <=  n_13910  AND n_13911;
inv_12364: n_13910  <= TRANSPORT NOT a_N2376  ;
delay_12365: n_13911  <= TRANSPORT a_SCH2ADDRREG_F5_G  ;
and1_12366: n_13912 <=  gnd;
delay_12367: a_LC1_F6  <= TRANSPORT a_EQ239  ;
xor2_12368: a_EQ239 <=  n_13915  XOR n_13922;
or2_12369: n_13915 <=  n_13916  OR n_13919;
and2_12370: n_13916 <=  n_13917  AND n_13918;
inv_12371: n_13917  <= TRANSPORT NOT a_N2377  ;
delay_12372: n_13918  <= TRANSPORT a_SCH3ADDRREG_F5_G  ;
and2_12373: n_13919 <=  n_13920  AND n_13921;
inv_12374: n_13920  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12375: n_13921  <= TRANSPORT a_SCH0ADDRREG_F5_G  ;
and1_12376: n_13922 <=  gnd;
dff_12377: DFF_a8237

    PORT MAP ( D => a_EQ039, CLK => a_LC3_F6_aCLK, CLRN => a_LC3_F6_aCLRN,
          PRN => vcc, Q => a_LC3_F6);
inv_12378: a_LC3_F6_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12379: a_EQ039 <=  n_13929  XOR n_13939;
or3_12380: n_13929 <=  n_13930  OR n_13933  OR n_13936;
and2_12381: n_13930 <=  n_13931  AND n_13932;
inv_12382: n_13931  <= TRANSPORT NOT startdma  ;
delay_12383: n_13932  <= TRANSPORT a_N423_aNOT  ;
and2_12384: n_13933 <=  n_13934  AND n_13935;
delay_12385: n_13934  <= TRANSPORT startdma  ;
delay_12386: n_13935  <= TRANSPORT a_LC2_F6  ;
and2_12387: n_13936 <=  n_13937  AND n_13938;
delay_12388: n_13937  <= TRANSPORT startdma  ;
delay_12389: n_13938  <= TRANSPORT a_LC1_F6  ;
and1_12390: n_13939 <=  gnd;
delay_12391: n_13940  <= TRANSPORT clk  ;
filter_12392: FILTER_a8237

    PORT MAP (IN1 => n_13940, Y => a_LC3_F6_aCLK);
delay_12393: a_N1726_aNOT  <= TRANSPORT a_EQ496  ;
xor2_12394: a_EQ496 <=  n_13944  XOR n_13951;
or2_12395: n_13944 <=  n_13945  OR n_13948;
and2_12396: n_13945 <=  n_13946  AND n_13947;
delay_12397: n_13946  <= TRANSPORT a_N2557  ;
delay_12398: n_13947  <= TRANSPORT a_N2546  ;
and2_12399: n_13948 <=  n_13949  AND n_13950;
inv_12400: n_13949  <= TRANSPORT NOT a_N2557  ;
delay_12401: n_13950  <= TRANSPORT a_LC4_F10  ;
and1_12402: n_13951 <=  gnd;
delay_12403: a_N1730  <= TRANSPORT a_EQ498  ;
xor2_12404: a_EQ498 <=  n_13954  XOR n_13961;
or2_12405: n_13954 <=  n_13955  OR n_13958;
and2_12406: n_13955 <=  n_13956  AND n_13957;
delay_12407: n_13956  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12408: n_13957  <= TRANSPORT a_SCH1ADDRREG_F6_G  ;
and2_12409: n_13958 <=  n_13959  AND n_13960;
inv_12410: n_13959  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12411: n_13960  <= TRANSPORT a_SCH0ADDRREG_F6_G  ;
and1_12412: n_13961 <=  gnd;
delay_12413: a_LC6_F10  <= TRANSPORT a_EQ492  ;
xor2_12414: a_EQ492 <=  n_13964  XOR n_13975;
or3_12415: n_13964 <=  n_13965  OR n_13968  OR n_13971;
and2_12416: n_13965 <=  n_13966  AND n_13967;
inv_12417: n_13966  <= TRANSPORT NOT a_N2557  ;
delay_12418: n_13967  <= TRANSPORT a_N1726_aNOT  ;
and2_12419: n_13968 <=  n_13969  AND n_13970;
inv_12420: n_13969  <= TRANSPORT NOT a_N2591  ;
delay_12421: n_13970  <= TRANSPORT a_N1726_aNOT  ;
and3_12422: n_13971 <=  n_13972  AND n_13973  AND n_13974;
delay_12423: n_13972  <= TRANSPORT a_N2557  ;
delay_12424: n_13973  <= TRANSPORT a_N2591  ;
delay_12425: n_13974  <= TRANSPORT a_N1730  ;
and1_12426: n_13975 <=  gnd;
delay_12427: a_LC2_F10  <= TRANSPORT a_EQ494  ;
xor2_12428: a_EQ494 <=  n_13978  XOR n_13985;
or2_12429: n_13978 <=  n_13979  OR n_13982;
and2_12430: n_13979 <=  n_13980  AND n_13981;
inv_12431: n_13980  <= TRANSPORT NOT a_N2376  ;
delay_12432: n_13981  <= TRANSPORT a_SCH2ADDRREG_F6_G  ;
and2_12433: n_13982 <=  n_13983  AND n_13984;
inv_12434: n_13983  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12435: n_13984  <= TRANSPORT a_SCH0ADDRREG_F6_G  ;
and1_12436: n_13985 <=  gnd;
delay_12437: a_LC3_F10  <= TRANSPORT a_EQ493  ;
xor2_12438: a_EQ493 <=  n_13988  XOR n_13995;
or2_12439: n_13988 <=  n_13989  OR n_13992;
and2_12440: n_13989 <=  n_13990  AND n_13991;
inv_12441: n_13990  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12442: n_13991  <= TRANSPORT a_SCH1ADDRREG_F6_G  ;
and2_12443: n_13992 <=  n_13993  AND n_13994;
inv_12444: n_13993  <= TRANSPORT NOT a_N2377  ;
delay_12445: n_13994  <= TRANSPORT a_SCH3ADDRREG_F6_G  ;
and1_12446: n_13995 <=  gnd;
dff_12447: DFF_a8237

    PORT MAP ( D => a_EQ038, CLK => a_LC4_F10_aCLK, CLRN => a_LC4_F10_aCLRN,
          PRN => vcc, Q => a_LC4_F10);
inv_12448: a_LC4_F10_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12449: a_EQ038 <=  n_14002  XOR n_14012;
or3_12450: n_14002 <=  n_14003  OR n_14006  OR n_14009;
and2_12451: n_14003 <=  n_14004  AND n_14005;
inv_12452: n_14004  <= TRANSPORT NOT startdma  ;
delay_12453: n_14005  <= TRANSPORT a_LC6_F10  ;
and2_12454: n_14006 <=  n_14007  AND n_14008;
delay_12455: n_14007  <= TRANSPORT startdma  ;
delay_12456: n_14008  <= TRANSPORT a_LC2_F10  ;
and2_12457: n_14009 <=  n_14010  AND n_14011;
delay_12458: n_14010  <= TRANSPORT startdma  ;
delay_12459: n_14011  <= TRANSPORT a_LC3_F10  ;
and1_12460: n_14012 <=  gnd;
delay_12461: n_14013  <= TRANSPORT clk  ;
filter_12462: FILTER_a8237

    PORT MAP (IN1 => n_14013, Y => a_LC4_F10_aCLK);
delay_12463: a_LC4_D27  <= TRANSPORT a_EQ200  ;
xor2_12464: a_EQ200 <=  n_14017  XOR n_14024;
or2_12465: n_14017 <=  n_14018  OR n_14021;
and2_12466: n_14018 <=  n_14019  AND n_14020;
delay_12467: n_14019  <= TRANSPORT a_N2557  ;
delay_12468: n_14020  <= TRANSPORT a_N2547  ;
and2_12469: n_14021 <=  n_14022  AND n_14023;
inv_12470: n_14022  <= TRANSPORT NOT a_N2557  ;
delay_12471: n_14023  <= TRANSPORT a_LC5_D27  ;
and1_12472: n_14024 <=  gnd;
delay_12473: a_LC3_D27  <= TRANSPORT a_EQ201  ;
xor2_12474: a_EQ201 <=  n_14027  XOR n_14034;
or2_12475: n_14027 <=  n_14028  OR n_14031;
and2_12476: n_14028 <=  n_14029  AND n_14030;
delay_12477: n_14029  <= TRANSPORT a_SNMEMR_aNOT  ;
delay_12478: n_14030  <= TRANSPORT a_SCH1ADDRREG_F7_G  ;
and2_12479: n_14031 <=  n_14032  AND n_14033;
inv_12480: n_14032  <= TRANSPORT NOT a_SNMEMR_aNOT  ;
delay_12481: n_14033  <= TRANSPORT a_SCH0ADDRREG_F7_G  ;
and1_12482: n_14034 <=  gnd;
delay_12483: a_N185_aNOT  <= TRANSPORT a_EQ205  ;
xor2_12484: a_EQ205 <=  n_14037  XOR n_14044;
or2_12485: n_14037 <=  n_14038  OR n_14041;
and2_12486: n_14038 <=  n_14039  AND n_14040;
inv_12487: n_14039  <= TRANSPORT NOT a_N2531  ;
delay_12488: n_14040  <= TRANSPORT a_LC4_D27  ;
and2_12489: n_14041 <=  n_14042  AND n_14043;
delay_12490: n_14042  <= TRANSPORT a_N2531  ;
delay_12491: n_14043  <= TRANSPORT a_LC3_D27  ;
and1_12492: n_14044 <=  gnd;
delay_12493: a_LC2_D27  <= TRANSPORT a_EQ203  ;
xor2_12494: a_EQ203 <=  n_14047  XOR n_14054;
or2_12495: n_14047 <=  n_14048  OR n_14051;
and2_12496: n_14048 <=  n_14049  AND n_14050;
inv_12497: n_14049  <= TRANSPORT NOT a_N2377  ;
delay_12498: n_14050  <= TRANSPORT a_SCH3ADDRREG_F7_G  ;
and2_12499: n_14051 <=  n_14052  AND n_14053;
inv_12500: n_14052  <= TRANSPORT NOT a_N2376  ;
delay_12501: n_14053  <= TRANSPORT a_SCH2ADDRREG_F7_G  ;
and1_12502: n_14054 <=  gnd;
delay_12503: a_LC1_D27  <= TRANSPORT a_EQ202  ;
xor2_12504: a_EQ202 <=  n_14057  XOR n_14064;
or2_12505: n_14057 <=  n_14058  OR n_14061;
and2_12506: n_14058 <=  n_14059  AND n_14060;
inv_12507: n_14059  <= TRANSPORT NOT a_N2598_aNOT  ;
delay_12508: n_14060  <= TRANSPORT a_SCH0ADDRREG_F7_G  ;
and2_12509: n_14061 <=  n_14062  AND n_14063;
inv_12510: n_14062  <= TRANSPORT NOT a_N88_aNOT  ;
delay_12511: n_14063  <= TRANSPORT a_SCH1ADDRREG_F7_G  ;
and1_12512: n_14064 <=  gnd;
dff_12513: DFF_a8237

    PORT MAP ( D => a_EQ037, CLK => a_LC5_D27_aCLK, CLRN => a_LC5_D27_aCLRN,
          PRN => vcc, Q => a_LC5_D27);
inv_12514: a_LC5_D27_aCLRN  <= TRANSPORT NOT reset  ;
xor2_12515: a_EQ037 <=  n_14071  XOR n_14081;
or3_12516: n_14071 <=  n_14072  OR n_14075  OR n_14078;
and2_12517: n_14072 <=  n_14073  AND n_14074;
inv_12518: n_14073  <= TRANSPORT NOT startdma  ;
delay_12519: n_14074  <= TRANSPORT a_N185_aNOT  ;
and2_12520: n_14075 <=  n_14076  AND n_14077;
delay_12521: n_14076  <= TRANSPORT startdma  ;
delay_12522: n_14077  <= TRANSPORT a_LC2_D27  ;
and2_12523: n_14078 <=  n_14079  AND n_14080;
delay_12524: n_14079  <= TRANSPORT startdma  ;
delay_12525: n_14080  <= TRANSPORT a_LC1_D27  ;
and1_12526: n_14081 <=  gnd;
delay_12527: n_14082  <= TRANSPORT clk  ;
filter_12528: FILTER_a8237

    PORT MAP (IN1 => n_14082, Y => a_LC5_D27_aCLK);
delay_12529: a_LC7_B10  <= TRANSPORT a_EQ110  ;
xor2_12530: a_EQ110 <=  n_14086  XOR n_14096;
or3_12531: n_14086 <=  n_14087  OR n_14090  OR n_14093;
and2_12532: n_14087 <=  n_14088  AND n_14089;
delay_12533: n_14088  <= TRANSPORT a_N1584  ;
delay_12534: n_14089  <= TRANSPORT a_STEMPORARYREG_F0_G  ;
and2_12535: n_14090 <=  n_14091  AND n_14092;
inv_12536: n_14091  <= TRANSPORT NOT a_N1584  ;
delay_12537: n_14092  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and2_12538: n_14093 <=  n_14094  AND n_14095;
inv_12539: n_14094  <= TRANSPORT NOT a_N2563_aNOT  ;
delay_12540: n_14095  <= TRANSPORT a_SADDRESSOUT_F8_G  ;
and1_12541: n_14096 <=  gnd;
delay_12542: a_SAEN_aNOT  <= TRANSPORT a_EQ864  ;
xor2_12543: a_EQ864 <=  n_14098  XOR n_14103;
or2_12544: n_14098 <=  n_14099  OR n_14101;
and1_12545: n_14099 <=  n_14100;
inv_12546: n_14100  <= TRANSPORT NOT a_N2563_aNOT  ;
and1_12547: n_14101 <=  n_14102;
inv_12548: n_14102  <= TRANSPORT NOT a_N1566  ;
and1_12549: n_14103 <=  gnd;
delay_12550: a_N2389  <= TRANSPORT a_EQ571  ;
xor2_12551: a_EQ571 <=  n_14106  XOR n_14111;
or2_12552: n_14106 <=  n_14107  OR n_14109;
and1_12553: n_14107 <=  n_14108;
delay_12554: n_14108  <= TRANSPORT a_N65  ;
and1_12555: n_14109 <=  n_14110;
inv_12556: n_14110  <= TRANSPORT NOT a_N75_aNOT  ;
and1_12557: n_14111 <=  gnd;
delay_12558: a_LC3_B9  <= TRANSPORT a_EQ121  ;
xor2_12559: a_EQ121 <=  n_14114  XOR n_14121;
or2_12560: n_14114 <=  n_14115  OR n_14118;
and2_12561: n_14115 <=  n_14116  AND n_14117;
inv_12562: n_14116  <= TRANSPORT NOT a_SMASKREG_F0_G_aNOT  ;
delay_12563: n_14117  <= TRANSPORT a_N2389  ;
and2_12564: n_14118 <=  n_14119  AND n_14120;
inv_12565: n_14119  <= TRANSPORT NOT a_N63_aNOT  ;
delay_12566: n_14120  <= TRANSPORT a_SREQUESTREG_F0_G  ;
and1_12567: n_14121 <=  gnd;
delay_12568: a_LC5_D23  <= TRANSPORT a_EQ111  ;
xor2_12569: a_EQ111 <=  n_14124  XOR n_14131;
or2_12570: n_14124 <=  n_14125  OR n_14128;
and2_12571: n_14125 <=  n_14126  AND n_14127;
inv_12572: n_14126  <= TRANSPORT NOT a_N77_aNOT  ;
delay_12573: n_14127  <= TRANSPORT a_SCH2ADDRREG_F8_G  ;
and2_12574: n_14128 <=  n_14129  AND n_14130;
inv_12575: n_14129  <= TRANSPORT NOT a_N2347  ;
delay_12576: n_14130  <= TRANSPORT a_SCH3WRDCNTREG_F8_G  ;
and1_12577: n_14131 <=  gnd;
delay_12578: a_LC2_F9  <= TRANSPORT a_EQ112  ;
xor2_12579: a_EQ112 <=  n_14134  XOR n_14141;
or2_12580: n_14134 <=  n_14135  OR n_14138;
and2_12581: n_14135 <=  n_14136  AND n_14137;
delay_12582: n_14136  <= TRANSPORT a_N2354_aNOT  ;
delay_12583: n_14137  <= TRANSPORT a_SCH0ADDRREG_F8_G  ;
and2_12584: n_14138 <=  n_14139  AND n_14140;
inv_12585: n_14139  <= TRANSPORT NOT a_N2348  ;
delay_12586: n_14140  <= TRANSPORT a_SCH3ADDRREG_F8_G  ;
and1_12587: n_14141 <=  gnd;
delay_12588: a_LC4_D23  <= TRANSPORT a_EQ113  ;
xor2_12589: a_EQ113 <=  n_14144  XOR n_14151;
or2_12590: n_14144 <=  n_14145  OR n_14148;
and2_12591: n_14145 <=  n_14146  AND n_14147;
inv_12592: n_14146  <= TRANSPORT NOT a_N2353  ;
delay_12593: n_14147  <= TRANSPORT a_SCH0WRDCNTREG_F8_G  ;
and2_12594: n_14148 <=  n_14149  AND n_14150;
inv_12595: n_14149  <= TRANSPORT NOT a_N2352  ;
delay_12596: n_14150  <= TRANSPORT a_SCH1ADDRREG_F8_G  ;
and1_12597: n_14151 <=  gnd;
delay_12598: a_LC3_D23  <= TRANSPORT a_EQ114  ;
xor2_12599: a_EQ114 <=  n_14154  XOR n_14162;
or2_12600: n_14154 <=  n_14155  OR n_14158;
and2_12601: n_14155 <=  n_14156  AND n_14157;
inv_12602: n_14156  <= TRANSPORT NOT a_N62_aNOT  ;
delay_12603: n_14157  <= TRANSPORT a_SCH2WRDCNTREG_F8_G  ;
and2_12604: n_14158 <=  n_14159  AND n_14161;
inv_12605: n_14159  <= TRANSPORT NOT a_N2351  ;
delay_12606: n_14161  <= TRANSPORT a_SCH1WRDCNTREG_F8_G  ;
and1_12607: n_14162 <=  gnd;
delay_12608: a_LC1_D23  <= TRANSPORT a_EQ115  ;
xor2_12609: a_EQ115 <=  n_14165  XOR n_14174;
or4_12610: n_14165 <=  n_14166  OR n_14168  OR n_14170  OR n_14172;
and1_12611: n_14166 <=  n_14167;
delay_12612: n_14167  <= TRANSPORT a_LC5_D23  ;
and1_12613: n_14168 <=  n_14169;
delay_12614: n_14169  <= TRANSPORT a_LC2_F9  ;
and1_12615: n_14170 <=  n_14171;
delay_12616: n_14171  <= TRANSPORT a_LC4_D23  ;
and1_12617: n_14172 <=  n_14173;
delay_12618: n_14173  <= TRANSPORT a_LC3_D23  ;
and1_12619: n_14174 <=  gnd;
delay_12620: a_LC6_D22  <= TRANSPORT a_EQ116  ;
xor2_12621: a_EQ116 <=  n_14177  XOR n_14184;
or2_12622: n_14177 <=  n_14178  OR n_14181;
and2_12623: n_14178 <=  n_14179  AND n_14180;
inv_12624: n_14179  <= TRANSPORT NOT a_N77_aNOT  ;
delay_12625: n_14180  <= TRANSPORT a_SCH2ADDRREG_F0_G  ;
and2_12626: n_14181 <=  n_14182  AND n_14183;
inv_12627: n_14182  <= TRANSPORT NOT a_N2347  ;
delay_12628: n_14183  <= TRANSPORT a_SCH3WRDCNTREG_F0_G  ;
and1_12629: n_14184 <=  gnd;
delay_12630: a_LC4_D22  <= TRANSPORT a_EQ117  ;
xor2_12631: a_EQ117 <=  n_14187  XOR n_14194;
or2_12632: n_14187 <=  n_14188  OR n_14191;
and2_12633: n_14188 <=  n_14189  AND n_14190;
delay_12634: n_14189  <= TRANSPORT a_N2354_aNOT  ;
delay_12635: n_14190  <= TRANSPORT a_SCH0ADDRREG_F0_G  ;
and2_12636: n_14191 <=  n_14192  AND n_14193;
inv_12637: n_14192  <= TRANSPORT NOT a_N2348  ;
delay_12638: n_14193  <= TRANSPORT a_SCH3ADDRREG_F0_G  ;
and1_12639: n_14194 <=  gnd;
delay_12640: a_LC2_D22  <= TRANSPORT a_EQ118  ;
xor2_12641: a_EQ118 <=  n_14197  XOR n_14204;
or2_12642: n_14197 <=  n_14198  OR n_14201;
and2_12643: n_14198 <=  n_14199  AND n_14200;
inv_12644: n_14199  <= TRANSPORT NOT a_N2353  ;
delay_12645: n_14200  <= TRANSPORT a_SCH0WRDCNTREG_F0_G  ;
and2_12646: n_14201 <=  n_14202  AND n_14203;
inv_12647: n_14202  <= TRANSPORT NOT a_N2352  ;
delay_12648: n_14203  <= TRANSPORT a_SCH1ADDRREG_F0_G  ;
and1_12649: n_14204 <=  gnd;
delay_12650: a_LC1_D22  <= TRANSPORT a_EQ119  ;
xor2_12651: a_EQ119 <=  n_14207  XOR n_14214;
or2_12652: n_14207 <=  n_14208  OR n_14211;
and2_12653: n_14208 <=  n_14209  AND n_14210;
inv_12654: n_14209  <= TRANSPORT NOT a_N62_aNOT  ;
delay_12655: n_14210  <= TRANSPORT a_SCH2WRDCNTREG_F0_G  ;
and2_12656: n_14211 <=  n_14212  AND n_14213;
inv_12657: n_14212  <= TRANSPORT NOT a_N2351  ;
delay_12658: n_14213  <= TRANSPORT a_SCH1WRDCNTREG_F0_G  ;
and1_12659: n_14214 <=  gnd;
delay_12660: a_LC5_D22  <= TRANSPORT a_EQ120  ;
xor2_12661: a_EQ120 <=  n_14217  XOR n_14226;
or4_12662: n_14217 <=  n_14218  OR n_14220  OR n_14222  OR n_14224;
and1_12663: n_14218 <=  n_14219;
delay_12664: n_14219  <= TRANSPORT a_LC6_D22  ;
and1_12665: n_14220 <=  n_14221;
delay_12666: n_14221  <= TRANSPORT a_LC4_D22  ;
and1_12667: n_14222 <=  n_14223;
delay_12668: n_14223  <= TRANSPORT a_LC2_D22  ;
and1_12669: n_14224 <=  n_14225;
delay_12670: n_14225  <= TRANSPORT a_LC1_D22  ;
and1_12671: n_14226 <=  gnd;
delay_12672: a_LC2_D23  <= TRANSPORT a_EQ122  ;
xor2_12673: a_EQ122 <=  n_14229  XOR n_14238;
or3_12674: n_14229 <=  n_14230  OR n_14232  OR n_14235;
and1_12675: n_14230 <=  n_14231;
delay_12676: n_14231  <= TRANSPORT a_LC3_B9  ;
and2_12677: n_14232 <=  n_14233  AND n_14234;
delay_12678: n_14233  <= TRANSPORT bytepointer  ;
delay_12679: n_14234  <= TRANSPORT a_LC1_D23  ;
and2_12680: n_14235 <=  n_14236  AND n_14237;
inv_12681: n_14236  <= TRANSPORT NOT bytepointer  ;
delay_12682: n_14237  <= TRANSPORT a_LC5_D22  ;
and1_12683: n_14238 <=  gnd;
delay_12684: a_N1830  <= TRANSPORT a_N1830_aIN  ;
xor2_12685: a_N1830_aIN <=  n_14241  XOR n_14244;
or1_12686: n_14241 <=  n_14242;
and1_12687: n_14242 <=  n_14243;
inv_12688: n_14243  <= TRANSPORT NOT a_LC4_A3  ;
and1_12689: n_14244 <=  gnd;
delay_12690: a_LC6_B10  <= TRANSPORT a_EQ123  ;
xor2_12691: a_EQ123 <=  n_14247  XOR n_14254;
or2_12692: n_14247 <=  n_14248  OR n_14251;
and2_12693: n_14248 <=  n_14249  AND n_14250;
delay_12694: n_14249  <= TRANSPORT a_STEMPORARYREG_F0_G  ;
delay_12695: n_14250  <= TRANSPORT a_N1830  ;
and2_12696: n_14251 <=  n_14252  AND n_14253;
inv_12697: n_14252  <= TRANSPORT NOT a_N2367  ;
delay_12698: n_14253  <= TRANSPORT a_STCSTATUS_F0_G  ;
and1_12699: n_14254 <=  gnd;
delay_12700: a_LC4_B10  <= TRANSPORT a_EQ124  ;
xor2_12701: a_EQ124 <=  n_14257  XOR n_14265;
or3_12702: n_14257 <=  n_14258  OR n_14260  OR n_14263;
and1_12703: n_14258 <=  n_14259;
delay_12704: n_14259  <= TRANSPORT a_LC6_B10  ;
and2_12705: n_14260 <=  n_14261  AND n_14262;
delay_12706: n_14261  <= TRANSPORT a_N73  ;
delay_12707: n_14262  <= TRANSPORT a_SCOMMANDREG_F0_G  ;
and1_12708: n_14263 <=  n_14264;
delay_12709: n_14264  <= TRANSPORT a_N66  ;
and1_12710: n_14265 <=  gnd;
delay_12711: a_G956  <= TRANSPORT a_EQ125  ;
xor2_12712: a_EQ125 <=  n_14267  XOR n_14277;
or3_12713: n_14267 <=  n_14268  OR n_14271  OR n_14274;
and2_12714: n_14268 <=  n_14269  AND n_14270;
delay_12715: n_14269  <= TRANSPORT a_LC7_B10  ;
inv_12716: n_14270  <= TRANSPORT NOT a_SAEN_aNOT  ;
and2_12717: n_14271 <=  n_14272  AND n_14273;
delay_12718: n_14272  <= TRANSPORT a_SAEN_aNOT  ;
delay_12719: n_14273  <= TRANSPORT a_LC2_D23  ;
and2_12720: n_14274 <=  n_14275  AND n_14276;
delay_12721: n_14275  <= TRANSPORT a_SAEN_aNOT  ;
delay_12722: n_14276  <= TRANSPORT a_LC4_B10  ;
and1_12723: n_14277 <=  gnd;
delay_12724: a_LC2_B21  <= TRANSPORT a_EQ143  ;
xor2_12725: a_EQ143 <=  n_14280  XOR n_14290;
or3_12726: n_14280 <=  n_14281  OR n_14284  OR n_14287;
and2_12727: n_14281 <=  n_14282  AND n_14283;
delay_12728: n_14282  <= TRANSPORT a_N1584  ;
delay_12729: n_14283  <= TRANSPORT a_STEMPORARYREG_F1_G  ;
and2_12730: n_14284 <=  n_14285  AND n_14286;
inv_12731: n_14285  <= TRANSPORT NOT a_N1584  ;
delay_12732: n_14286  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
and2_12733: n_14287 <=  n_14288  AND n_14289;
inv_12734: n_14288  <= TRANSPORT NOT a_N2563_aNOT  ;
delay_12735: n_14289  <= TRANSPORT a_SADDRESSOUT_F9_G  ;
and1_12736: n_14290 <=  gnd;
delay_12737: a_LC8_C8  <= TRANSPORT a_EQ152  ;
xor2_12738: a_EQ152 <=  n_14293  XOR n_14300;
or2_12739: n_14293 <=  n_14294  OR n_14297;
and2_12740: n_14294 <=  n_14295  AND n_14296;
inv_12741: n_14295  <= TRANSPORT NOT a_N2352  ;
delay_12742: n_14296  <= TRANSPORT a_SCH1ADDRREG_F1_G  ;
and2_12743: n_14297 <=  n_14298  AND n_14299;
inv_12744: n_14298  <= TRANSPORT NOT a_N2347  ;
delay_12745: n_14299  <= TRANSPORT a_SCH3WRDCNTREG_F1_G  ;
and1_12746: n_14300 <=  gnd;
delay_12747: a_LC7_C8  <= TRANSPORT a_EQ153  ;
xor2_12748: a_EQ153 <=  n_14303  XOR n_14310;
or2_12749: n_14303 <=  n_14304  OR n_14307;
and2_12750: n_14304 <=  n_14305  AND n_14306;
inv_12751: n_14305  <= TRANSPORT NOT a_N2353  ;
delay_12752: n_14306  <= TRANSPORT a_SCH0WRDCNTREG_F1_G  ;
and2_12753: n_14307 <=  n_14308  AND n_14309;
inv_12754: n_14308  <= TRANSPORT NOT a_N2351  ;
delay_12755: n_14309  <= TRANSPORT a_SCH1WRDCNTREG_F1_G  ;
and1_12756: n_14310 <=  gnd;
delay_12757: a_LC5_C8  <= TRANSPORT a_EQ154  ;
xor2_12758: a_EQ154 <=  n_14313  XOR n_14320;
or2_12759: n_14313 <=  n_14314  OR n_14317;
and2_12760: n_14314 <=  n_14315  AND n_14316;
inv_12761: n_14315  <= TRANSPORT NOT a_N77_aNOT  ;
delay_12762: n_14316  <= TRANSPORT a_SCH2ADDRREG_F1_G  ;
and2_12763: n_14317 <=  n_14318  AND n_14319;
delay_12764: n_14318  <= TRANSPORT a_N2354_aNOT  ;
delay_12765: n_14319  <= TRANSPORT a_SCH0ADDRREG_F1_G  ;
and1_12766: n_14320 <=  gnd;
delay_12767: a_LC4_C8  <= TRANSPORT a_EQ155  ;
xor2_12768: a_EQ155 <=  n_14323  XOR n_14330;
or2_12769: n_14323 <=  n_14324  OR n_14327;
and2_12770: n_14324 <=  n_14325  AND n_14326;
inv_12771: n_14325  <= TRANSPORT NOT a_N62_aNOT  ;
delay_12772: n_14326  <= TRANSPORT a_SCH2WRDCNTREG_F1_G  ;
and2_12773: n_14327 <=  n_14328  AND n_14329;
inv_12774: n_14328  <= TRANSPORT NOT a_N2348  ;
delay_12775: n_14329  <= TRANSPORT a_SCH3ADDRREG_F1_G  ;
and1_12776: n_14330 <=  gnd;
delay_12777: a_LC6_C8  <= TRANSPORT a_EQ156  ;
xor2_12778: a_EQ156 <=  n_14333  XOR n_14342;
or4_12779: n_14333 <=  n_14334  OR n_14336  OR n_14338  OR n_14340;
and1_12780: n_14334 <=  n_14335;
delay_12781: n_14335  <= TRANSPORT a_LC8_C8  ;
and1_12782: n_14336 <=  n_14337;
delay_12783: n_14337  <= TRANSPORT a_LC7_C8  ;
and1_12784: n_14338 <=  n_14339;
delay_12785: n_14339  <= TRANSPORT a_LC5_C8  ;
and1_12786: n_14340 <=  n_14341;
delay_12787: n_14341  <= TRANSPORT a_LC4_C8  ;
and1_12788: n_14342 <=  gnd;
delay_12789: a_LC4_A17  <= TRANSPORT a_EQ148  ;
xor2_12790: a_EQ148 <=  n_14345  XOR n_14352;
or2_12791: n_14345 <=  n_14346  OR n_14349;
and2_12792: n_14346 <=  n_14347  AND n_14348;
inv_12793: n_14347  <= TRANSPORT NOT a_N2353  ;
delay_12794: n_14348  <= TRANSPORT a_SCH0WRDCNTREG_F9_G  ;
and2_12795: n_14349 <=  n_14350  AND n_14351;
inv_12796: n_14350  <= TRANSPORT NOT a_N2351  ;
delay_12797: n_14351  <= TRANSPORT a_SCH1WRDCNTREG_F9_G  ;
and1_12798: n_14352 <=  gnd;
delay_12799: a_LC3_A17  <= TRANSPORT a_EQ149  ;
xor2_12800: a_EQ149 <=  n_14355  XOR n_14362;
or2_12801: n_14355 <=  n_14356  OR n_14359;
and2_12802: n_14356 <=  n_14357  AND n_14358;
inv_12803: n_14357  <= TRANSPORT NOT a_N77_aNOT  ;
delay_12804: n_14358  <= TRANSPORT a_SCH2ADDRREG_F9_G  ;
and2_12805: n_14359 <=  n_14360  AND n_14361;
delay_12806: n_14360  <= TRANSPORT a_N2354_aNOT  ;
delay_12807: n_14361  <= TRANSPORT a_SCH0ADDRREG_F9_G  ;
and1_12808: n_14362 <=  gnd;
delay_12809: a_LC2_A17  <= TRANSPORT a_EQ150  ;
xor2_12810: a_EQ150 <=  n_14365  XOR n_14372;
or2_12811: n_14365 <=  n_14366  OR n_14369;
and2_12812: n_14366 <=  n_14367  AND n_14368;
inv_12813: n_14367  <= TRANSPORT NOT a_N62_aNOT  ;
delay_12814: n_14368  <= TRANSPORT a_SCH2WRDCNTREG_F9_G  ;
and2_12815: n_14369 <=  n_14370  AND n_14371;
inv_12816: n_14370  <= TRANSPORT NOT a_N2348  ;
delay_12817: n_14371  <= TRANSPORT a_SCH3ADDRREG_F9_G  ;
and1_12818: n_14372 <=  gnd;
delay_12819: a_LC1_A17  <= TRANSPORT a_EQ151  ;
xor2_12820: a_EQ151 <=  n_14375  XOR n_14382;
or3_12821: n_14375 <=  n_14376  OR n_14378  OR n_14380;
and1_12822: n_14376 <=  n_14377;
delay_12823: n_14377  <= TRANSPORT a_LC4_A17  ;
and1_12824: n_14378 <=  n_14379;
delay_12825: n_14379  <= TRANSPORT a_LC3_A17  ;
and1_12826: n_14380 <=  n_14381;
delay_12827: n_14381  <= TRANSPORT a_LC2_A17  ;
and1_12828: n_14382 <=  gnd;
delay_12829: a_LC5_A17  <= TRANSPORT a_EQ147  ;
xor2_12830: a_EQ147 <=  n_14385  XOR n_14392;
or2_12831: n_14385 <=  n_14386  OR n_14389;
and2_12832: n_14386 <=  n_14387  AND n_14388;
inv_12833: n_14387  <= TRANSPORT NOT a_N2352  ;
delay_12834: n_14388  <= TRANSPORT a_SCH1ADDRREG_F9_G  ;
and2_12835: n_14389 <=  n_14390  AND n_14391;
inv_12836: n_14390  <= TRANSPORT NOT a_N2347  ;
delay_12837: n_14391  <= TRANSPORT a_SCH3WRDCNTREG_F9_G  ;
and1_12838: n_14392 <=  gnd;
delay_12839: a_LC6_A17  <= TRANSPORT a_EQ157  ;
xor2_12840: a_EQ157 <=  n_14395  XOR n_14405;
or3_12841: n_14395 <=  n_14396  OR n_14399  OR n_14402;
and2_12842: n_14396 <=  n_14397  AND n_14398;
inv_12843: n_14397  <= TRANSPORT NOT bytepointer  ;
delay_12844: n_14398  <= TRANSPORT a_LC6_C8  ;
and2_12845: n_14399 <=  n_14400  AND n_14401;
delay_12846: n_14400  <= TRANSPORT bytepointer  ;
delay_12847: n_14401  <= TRANSPORT a_LC1_A17  ;
and2_12848: n_14402 <=  n_14403  AND n_14404;
delay_12849: n_14403  <= TRANSPORT bytepointer  ;
delay_12850: n_14404  <= TRANSPORT a_LC5_A17  ;
and1_12851: n_14405 <=  gnd;
delay_12852: a_LC5_B23  <= TRANSPORT a_EQ145  ;
xor2_12853: a_EQ145 <=  n_14408  XOR n_14415;
or2_12854: n_14408 <=  n_14409  OR n_14412;
and2_12855: n_14409 <=  n_14410  AND n_14411;
inv_12856: n_14410  <= TRANSPORT NOT a_N63_aNOT  ;
delay_12857: n_14411  <= TRANSPORT a_SREQUESTREG_F1_G  ;
and2_12858: n_14412 <=  n_14413  AND n_14414;
inv_12859: n_14413  <= TRANSPORT NOT a_N2367  ;
delay_12860: n_14414  <= TRANSPORT a_STCSTATUS_F1_G  ;
and1_12861: n_14415 <=  gnd;
delay_12862: a_LC5_B21  <= TRANSPORT a_EQ146  ;
xor2_12863: a_EQ146 <=  n_14418  XOR n_14426;
or3_12864: n_14418 <=  n_14419  OR n_14421  OR n_14424;
and1_12865: n_14419 <=  n_14420;
delay_12866: n_14420  <= TRANSPORT a_LC5_B23  ;
and2_12867: n_14421 <=  n_14422  AND n_14423;
inv_12868: n_14422  <= TRANSPORT NOT a_LC4_A3  ;
delay_12869: n_14423  <= TRANSPORT a_STEMPORARYREG_F1_G  ;
and1_12870: n_14424 <=  n_14425;
delay_12871: n_14425  <= TRANSPORT a_N66  ;
and1_12872: n_14426 <=  gnd;
delay_12873: a_LC4_B21  <= TRANSPORT a_EQ144  ;
xor2_12874: a_EQ144 <=  n_14429  XOR n_14436;
or2_12875: n_14429 <=  n_14430  OR n_14433;
and2_12876: n_14430 <=  n_14431  AND n_14432;
inv_12877: n_14431  <= TRANSPORT NOT a_SMASKREG_F1_G_aNOT  ;
delay_12878: n_14432  <= TRANSPORT a_N2389  ;
and2_12879: n_14433 <=  n_14434  AND n_14435;
delay_12880: n_14434  <= TRANSPORT a_N73  ;
delay_12881: n_14435  <= TRANSPORT a_SCOMMANDREG_F1_G  ;
and1_12882: n_14436 <=  gnd;
delay_12883: a_LC7_B21  <= TRANSPORT a_EQ158  ;
xor2_12884: a_EQ158 <=  n_14439  XOR n_14446;
or3_12885: n_14439 <=  n_14440  OR n_14442  OR n_14444;
and1_12886: n_14440 <=  n_14441;
delay_12887: n_14441  <= TRANSPORT a_LC6_A17  ;
and1_12888: n_14442 <=  n_14443;
delay_12889: n_14443  <= TRANSPORT a_LC5_B21  ;
and1_12890: n_14444 <=  n_14445;
delay_12891: n_14445  <= TRANSPORT a_LC4_B21  ;
and1_12892: n_14446 <=  gnd;
delay_12893: a_G1027  <= TRANSPORT a_EQ159  ;
xor2_12894: a_EQ159 <=  n_14448  XOR n_14459;
or3_12895: n_14448 <=  n_14449  OR n_14453  OR n_14456;
and3_12896: n_14449 <=  n_14450  AND n_14451  AND n_14452;
delay_12897: n_14450  <= TRANSPORT a_N2563_aNOT  ;
delay_12898: n_14451  <= TRANSPORT a_N1566  ;
delay_12899: n_14452  <= TRANSPORT a_LC2_B21  ;
and2_12900: n_14453 <=  n_14454  AND n_14455;
inv_12901: n_14454  <= TRANSPORT NOT a_N2563_aNOT  ;
delay_12902: n_14455  <= TRANSPORT a_LC7_B21  ;
and2_12903: n_14456 <=  n_14457  AND n_14458;
inv_12904: n_14457  <= TRANSPORT NOT a_N1566  ;
delay_12905: n_14458  <= TRANSPORT a_LC7_B21  ;
and1_12906: n_14459 <=  gnd;
delay_12907: a_LC7_E23  <= TRANSPORT a_EQ077  ;
xor2_12908: a_EQ077 <=  n_14462  XOR n_14472;
or3_12909: n_14462 <=  n_14463  OR n_14466  OR n_14469;
and2_12910: n_14463 <=  n_14464  AND n_14465;
delay_12911: n_14464  <= TRANSPORT a_N1584  ;
delay_12912: n_14465  <= TRANSPORT a_STEMPORARYREG_F2_G  ;
and2_12913: n_14466 <=  n_14467  AND n_14468;
inv_12914: n_14467  <= TRANSPORT NOT a_N1584  ;
delay_12915: n_14468  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and2_12916: n_14469 <=  n_14470  AND n_14471;
inv_12917: n_14470  <= TRANSPORT NOT a_N2563_aNOT  ;
delay_12918: n_14471  <= TRANSPORT a_SADDRESSOUT_F10_G  ;
and1_12919: n_14472 <=  gnd;
delay_12920: a_LC8_E26  <= TRANSPORT a_EQ480  ;
xor2_12921: a_EQ480 <=  n_14475  XOR n_14484;
or2_12922: n_14475 <=  n_14476  OR n_14480;
and3_12923: n_14476 <=  n_14477  AND n_14478  AND n_14479;
inv_12924: n_14477  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
inv_12925: n_14478  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_12926: n_14479  <= TRANSPORT a_SCH0MODEREG_F0_G  ;
and3_12927: n_14480 <=  n_14481  AND n_14482  AND n_14483;
delay_12928: n_14481  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_12929: n_14482  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_12930: n_14483  <= TRANSPORT a_SCH2MODEREG_F0_G  ;
and1_12931: n_14484 <=  gnd;
delay_12932: a_LC7_E26  <= TRANSPORT a_EQ481  ;
xor2_12933: a_EQ481 <=  n_14487  XOR n_14496;
or2_12934: n_14487 <=  n_14488  OR n_14492;
and3_12935: n_14488 <=  n_14489  AND n_14490  AND n_14491;
delay_12936: n_14489  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
delay_12937: n_14490  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
delay_12938: n_14491  <= TRANSPORT a_SCH3MODEREG_F0_G  ;
and3_12939: n_14492 <=  n_14493  AND n_14494  AND n_14495;
inv_12940: n_14493  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_12941: n_14494  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
delay_12942: n_14495  <= TRANSPORT a_SCH1MODEREG_F0_G  ;
and1_12943: n_14496 <=  gnd;
delay_12944: a_N1647_aNOT  <= TRANSPORT a_EQ482  ;
xor2_12945: a_EQ482 <=  n_14499  XOR n_14506;
or2_12946: n_14499 <=  n_14500  OR n_14503;
and2_12947: n_14500 <=  n_14501  AND n_14502;
delay_12948: n_14501  <= TRANSPORT a_N66  ;
delay_12949: n_14502  <= TRANSPORT a_LC8_E26  ;
and2_12950: n_14503 <=  n_14504  AND n_14505;
delay_12951: n_14504  <= TRANSPORT a_N66  ;
delay_12952: n_14505  <= TRANSPORT a_LC7_E26  ;
and1_12953: n_14506 <=  gnd;
delay_12954: a_LC6_B7  <= TRANSPORT a_EQ090  ;
xor2_12955: a_EQ090 <=  n_14509  XOR n_14516;
or2_12956: n_14509 <=  n_14510  OR n_14513;
and2_12957: n_14510 <=  n_14511  AND n_14512;
inv_12958: n_14511  <= TRANSPORT NOT a_N63_aNOT  ;
delay_12959: n_14512  <= TRANSPORT a_SREQUESTREG_F2_G  ;
and2_12960: n_14513 <=  n_14514  AND n_14515;
inv_12961: n_14514  <= TRANSPORT NOT a_N2367  ;
delay_12962: n_14515  <= TRANSPORT a_STCSTATUS_F2_G  ;
and1_12963: n_14516 <=  gnd;
delay_12964: a_LC8_E23  <= TRANSPORT a_EQ091  ;
xor2_12965: a_EQ091 <=  n_14519  XOR n_14527;
or3_12966: n_14519 <=  n_14520  OR n_14522  OR n_14524;
and1_12967: n_14520 <=  n_14521;
delay_12968: n_14521  <= TRANSPORT a_N1647_aNOT  ;
and1_12969: n_14522 <=  n_14523;
delay_12970: n_14523  <= TRANSPORT a_LC6_B7  ;
and2_12971: n_14524 <=  n_14525  AND n_14526;
inv_12972: n_14525  <= TRANSPORT NOT a_LC4_A3  ;
delay_12973: n_14526  <= TRANSPORT a_STEMPORARYREG_F2_G  ;
and1_12974: n_14527 <=  gnd;
delay_12975: a_LC4_B14  <= TRANSPORT a_EQ088  ;
xor2_12976: a_EQ088 <=  n_14530  XOR n_14537;
or2_12977: n_14530 <=  n_14531  OR n_14534;
and2_12978: n_14531 <=  n_14532  AND n_14533;
inv_12979: n_14532  <= TRANSPORT NOT a_SMASKREG_F2_G_aNOT  ;
delay_12980: n_14533  <= TRANSPORT a_N2389  ;
and2_12981: n_14534 <=  n_14535  AND n_14536;
delay_12982: n_14535  <= TRANSPORT a_N73  ;
delay_12983: n_14536  <= TRANSPORT a_SCOMMANDREG_F2_G  ;
and1_12984: n_14537 <=  gnd;
delay_12985: a_LC2_C21  <= TRANSPORT a_EQ078  ;
xor2_12986: a_EQ078 <=  n_14540  XOR n_14547;
or2_12987: n_14540 <=  n_14541  OR n_14544;
and2_12988: n_14541 <=  n_14542  AND n_14543;
inv_12989: n_14542  <= TRANSPORT NOT a_N77_aNOT  ;
delay_12990: n_14543  <= TRANSPORT a_SCH2ADDRREG_F2_G  ;
and2_12991: n_14544 <=  n_14545  AND n_14546;
inv_12992: n_14545  <= TRANSPORT NOT a_N2347  ;
delay_12993: n_14546  <= TRANSPORT a_SCH3WRDCNTREG_F2_G  ;
and1_12994: n_14547 <=  gnd;
delay_12995: a_LC7_C21  <= TRANSPORT a_EQ079  ;
xor2_12996: a_EQ079 <=  n_14550  XOR n_14557;
or2_12997: n_14550 <=  n_14551  OR n_14554;
and2_12998: n_14551 <=  n_14552  AND n_14553;
inv_12999: n_14552  <= TRANSPORT NOT a_N2348  ;
delay_13000: n_14553  <= TRANSPORT a_SCH3ADDRREG_F2_G  ;
and2_13001: n_14554 <=  n_14555  AND n_14556;
inv_13002: n_14555  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13003: n_14556  <= TRANSPORT a_SCH2WRDCNTREG_F2_G  ;
and1_13004: n_14557 <=  gnd;
delay_13005: a_LC6_C21  <= TRANSPORT a_EQ080  ;
xor2_13006: a_EQ080 <=  n_14560  XOR n_14567;
or2_13007: n_14560 <=  n_14561  OR n_14564;
and2_13008: n_14561 <=  n_14562  AND n_14563;
inv_13009: n_14562  <= TRANSPORT NOT a_N2352  ;
delay_13010: n_14563  <= TRANSPORT a_SCH1ADDRREG_F2_G  ;
and2_13011: n_14564 <=  n_14565  AND n_14566;
inv_13012: n_14565  <= TRANSPORT NOT a_N2353  ;
delay_13013: n_14566  <= TRANSPORT a_SCH0WRDCNTREG_F2_G  ;
and1_13014: n_14567 <=  gnd;
delay_13015: a_LC4_C21  <= TRANSPORT a_EQ081  ;
xor2_13016: a_EQ081 <=  n_14570  XOR n_14577;
or2_13017: n_14570 <=  n_14571  OR n_14574;
and2_13018: n_14571 <=  n_14572  AND n_14573;
delay_13019: n_14572  <= TRANSPORT a_N2354_aNOT  ;
delay_13020: n_14573  <= TRANSPORT a_SCH0ADDRREG_F2_G  ;
and2_13021: n_14574 <=  n_14575  AND n_14576;
inv_13022: n_14575  <= TRANSPORT NOT a_N2351  ;
delay_13023: n_14576  <= TRANSPORT a_SCH1WRDCNTREG_F2_G  ;
and1_13024: n_14577 <=  gnd;
delay_13025: a_LC5_C21  <= TRANSPORT a_EQ082  ;
xor2_13026: a_EQ082 <=  n_14580  XOR n_14589;
or4_13027: n_14580 <=  n_14581  OR n_14583  OR n_14585  OR n_14587;
and1_13028: n_14581 <=  n_14582;
delay_13029: n_14582  <= TRANSPORT a_LC2_C21  ;
and1_13030: n_14583 <=  n_14584;
delay_13031: n_14584  <= TRANSPORT a_LC7_C21  ;
and1_13032: n_14585 <=  n_14586;
delay_13033: n_14586  <= TRANSPORT a_LC6_C21  ;
and1_13034: n_14587 <=  n_14588;
delay_13035: n_14588  <= TRANSPORT a_LC4_C21  ;
and1_13036: n_14589 <=  gnd;
delay_13037: a_LC5_E4  <= TRANSPORT a_EQ083  ;
xor2_13038: a_EQ083 <=  n_14592  XOR n_14599;
or2_13039: n_14592 <=  n_14593  OR n_14596;
and2_13040: n_14593 <=  n_14594  AND n_14595;
inv_13041: n_14594  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13042: n_14595  <= TRANSPORT a_SCH2ADDRREG_F10_G  ;
and2_13043: n_14596 <=  n_14597  AND n_14598;
inv_13044: n_14597  <= TRANSPORT NOT a_N2347  ;
delay_13045: n_14598  <= TRANSPORT a_SH3WRDCNTREG_F10_G  ;
and1_13046: n_14599 <=  gnd;
delay_13047: a_LC4_E4  <= TRANSPORT a_EQ084  ;
xor2_13048: a_EQ084 <=  n_14602  XOR n_14609;
or2_13049: n_14602 <=  n_14603  OR n_14606;
and2_13050: n_14603 <=  n_14604  AND n_14605;
inv_13051: n_14604  <= TRANSPORT NOT a_N2348  ;
delay_13052: n_14605  <= TRANSPORT a_SCH3ADDRREG_F10_G  ;
and2_13053: n_14606 <=  n_14607  AND n_14608;
inv_13054: n_14607  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13055: n_14608  <= TRANSPORT a_SH2WRDCNTREG_F10_G  ;
and1_13056: n_14609 <=  gnd;
delay_13057: a_LC4_E27  <= TRANSPORT a_EQ085  ;
xor2_13058: a_EQ085 <=  n_14612  XOR n_14619;
or2_13059: n_14612 <=  n_14613  OR n_14616;
and2_13060: n_14613 <=  n_14614  AND n_14615;
inv_13061: n_14614  <= TRANSPORT NOT a_N2352  ;
delay_13062: n_14615  <= TRANSPORT a_SCH1ADDRREG_F10_G  ;
and2_13063: n_14616 <=  n_14617  AND n_14618;
inv_13064: n_14617  <= TRANSPORT NOT a_N2353  ;
delay_13065: n_14618  <= TRANSPORT a_SH0WRDCNTREG_F10_G  ;
and1_13066: n_14619 <=  gnd;
delay_13067: a_LC2_E18  <= TRANSPORT a_EQ086  ;
xor2_13068: a_EQ086 <=  n_14622  XOR n_14629;
or2_13069: n_14622 <=  n_14623  OR n_14626;
and2_13070: n_14623 <=  n_14624  AND n_14625;
delay_13071: n_14624  <= TRANSPORT a_N2354_aNOT  ;
delay_13072: n_14625  <= TRANSPORT a_SCH0ADDRREG_F10_G  ;
and2_13073: n_14626 <=  n_14627  AND n_14628;
inv_13074: n_14627  <= TRANSPORT NOT a_N2351  ;
delay_13075: n_14628  <= TRANSPORT a_SH1WRDCNTREG_F10_G  ;
and1_13076: n_14629 <=  gnd;
delay_13077: a_LC3_E4  <= TRANSPORT a_EQ087  ;
xor2_13078: a_EQ087 <=  n_14632  XOR n_14641;
or4_13079: n_14632 <=  n_14633  OR n_14635  OR n_14637  OR n_14639;
and1_13080: n_14633 <=  n_14634;
delay_13081: n_14634  <= TRANSPORT a_LC5_E4  ;
and1_13082: n_14635 <=  n_14636;
delay_13083: n_14636  <= TRANSPORT a_LC4_E4  ;
and1_13084: n_14637 <=  n_14638;
delay_13085: n_14638  <= TRANSPORT a_LC4_E27  ;
and1_13086: n_14639 <=  n_14640;
delay_13087: n_14640  <= TRANSPORT a_LC2_E18  ;
and1_13088: n_14641 <=  gnd;
delay_13089: a_LC6_E4  <= TRANSPORT a_EQ089  ;
xor2_13090: a_EQ089 <=  n_14644  XOR n_14653;
or3_13091: n_14644 <=  n_14645  OR n_14647  OR n_14650;
and1_13092: n_14645 <=  n_14646;
delay_13093: n_14646  <= TRANSPORT a_LC4_B14  ;
and2_13094: n_14647 <=  n_14648  AND n_14649;
inv_13095: n_14648  <= TRANSPORT NOT bytepointer  ;
delay_13096: n_14649  <= TRANSPORT a_LC5_C21  ;
and2_13097: n_14650 <=  n_14651  AND n_14652;
delay_13098: n_14651  <= TRANSPORT bytepointer  ;
delay_13099: n_14652  <= TRANSPORT a_LC3_E4  ;
and1_13100: n_14653 <=  gnd;
delay_13101: a_G200  <= TRANSPORT a_EQ092  ;
xor2_13102: a_EQ092 <=  n_14655  XOR n_14665;
or3_13103: n_14655 <=  n_14656  OR n_14659  OR n_14662;
and2_13104: n_14656 <=  n_14657  AND n_14658;
inv_13105: n_14657  <= TRANSPORT NOT a_SAEN_aNOT  ;
delay_13106: n_14658  <= TRANSPORT a_LC7_E23  ;
and2_13107: n_14659 <=  n_14660  AND n_14661;
delay_13108: n_14660  <= TRANSPORT a_SAEN_aNOT  ;
delay_13109: n_14661  <= TRANSPORT a_LC8_E23  ;
and2_13110: n_14662 <=  n_14663  AND n_14664;
delay_13111: n_14663  <= TRANSPORT a_SAEN_aNOT  ;
delay_13112: n_14664  <= TRANSPORT a_LC6_E4  ;
and1_13113: n_14665 <=  gnd;
delay_13114: a_LC2_A27  <= TRANSPORT a_EQ060  ;
xor2_13115: a_EQ060 <=  n_14668  XOR n_14675;
or2_13116: n_14668 <=  n_14669  OR n_14672;
and2_13117: n_14669 <=  n_14670  AND n_14671;
delay_13118: n_14670  <= TRANSPORT a_N1584  ;
delay_13119: n_14671  <= TRANSPORT a_STEMPORARYREG_F3_G  ;
and2_13120: n_14672 <=  n_14673  AND n_14674;
inv_13121: n_14673  <= TRANSPORT NOT a_N1584  ;
delay_13122: n_14674  <= TRANSPORT a_SADDRESSOUT_F11_G  ;
and1_13123: n_14675 <=  gnd;
delay_13124: a_LC6_A10  <= TRANSPORT a_EQ066  ;
xor2_13125: a_EQ066 <=  n_14678  XOR n_14685;
or2_13126: n_14678 <=  n_14679  OR n_14682;
and2_13127: n_14679 <=  n_14680  AND n_14681;
delay_13128: n_14680  <= TRANSPORT a_N2354_aNOT  ;
delay_13129: n_14681  <= TRANSPORT a_SCH0ADDRREG_F11_G  ;
and2_13130: n_14682 <=  n_14683  AND n_14684;
inv_13131: n_14683  <= TRANSPORT NOT a_N2347  ;
delay_13132: n_14684  <= TRANSPORT a_SH3WRDCNTREG_F11_G  ;
and1_13133: n_14685 <=  gnd;
delay_13134: a_LC5_A10  <= TRANSPORT a_EQ067  ;
xor2_13135: a_EQ067 <=  n_14688  XOR n_14695;
or2_13136: n_14688 <=  n_14689  OR n_14692;
and2_13137: n_14689 <=  n_14690  AND n_14691;
inv_13138: n_14690  <= TRANSPORT NOT a_N2353  ;
delay_13139: n_14691  <= TRANSPORT a_SH0WRDCNTREG_F11_G  ;
and2_13140: n_14692 <=  n_14693  AND n_14694;
inv_13141: n_14693  <= TRANSPORT NOT a_N2352  ;
delay_13142: n_14694  <= TRANSPORT a_SCH1ADDRREG_F11_G  ;
and1_13143: n_14695 <=  gnd;
delay_13144: a_LC4_A10  <= TRANSPORT a_EQ068  ;
xor2_13145: a_EQ068 <=  n_14698  XOR n_14705;
or2_13146: n_14698 <=  n_14699  OR n_14702;
and2_13147: n_14699 <=  n_14700  AND n_14701;
inv_13148: n_14700  <= TRANSPORT NOT a_N2348  ;
delay_13149: n_14701  <= TRANSPORT a_SCH3ADDRREG_F11_G  ;
and2_13150: n_14702 <=  n_14703  AND n_14704;
inv_13151: n_14703  <= TRANSPORT NOT a_N2351  ;
delay_13152: n_14704  <= TRANSPORT a_SH1WRDCNTREG_F11_G  ;
and1_13153: n_14705 <=  gnd;
delay_13154: a_LC3_A10  <= TRANSPORT a_EQ069  ;
xor2_13155: a_EQ069 <=  n_14708  XOR n_14715;
or2_13156: n_14708 <=  n_14709  OR n_14712;
and2_13157: n_14709 <=  n_14710  AND n_14711;
inv_13158: n_14710  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13159: n_14711  <= TRANSPORT a_SCH2ADDRREG_F11_G  ;
and2_13160: n_14712 <=  n_14713  AND n_14714;
inv_13161: n_14713  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13162: n_14714  <= TRANSPORT a_SH2WRDCNTREG_F11_G  ;
and1_13163: n_14715 <=  gnd;
delay_13164: a_LC1_A10  <= TRANSPORT a_EQ070  ;
xor2_13165: a_EQ070 <=  n_14718  XOR n_14727;
or4_13166: n_14718 <=  n_14719  OR n_14721  OR n_14723  OR n_14725;
and1_13167: n_14719 <=  n_14720;
delay_13168: n_14720  <= TRANSPORT a_LC6_A10  ;
and1_13169: n_14721 <=  n_14722;
delay_13170: n_14722  <= TRANSPORT a_LC5_A10  ;
and1_13171: n_14723 <=  n_14724;
delay_13172: n_14724  <= TRANSPORT a_LC4_A10  ;
and1_13173: n_14725 <=  n_14726;
delay_13174: n_14726  <= TRANSPORT a_LC3_A10  ;
and1_13175: n_14727 <=  gnd;
delay_13176: a_LC6_C13  <= TRANSPORT a_EQ062  ;
xor2_13177: a_EQ062 <=  n_14730  XOR n_14737;
or2_13178: n_14730 <=  n_14731  OR n_14734;
and2_13179: n_14731 <=  n_14732  AND n_14733;
inv_13180: n_14732  <= TRANSPORT NOT a_N2353  ;
delay_13181: n_14733  <= TRANSPORT a_SCH0WRDCNTREG_F3_G  ;
and2_13182: n_14734 <=  n_14735  AND n_14736;
inv_13183: n_14735  <= TRANSPORT NOT a_N2352  ;
delay_13184: n_14736  <= TRANSPORT a_SCH1ADDRREG_F3_G  ;
and1_13185: n_14737 <=  gnd;
delay_13186: a_LC3_C8  <= TRANSPORT a_EQ063  ;
xor2_13187: a_EQ063 <=  n_14740  XOR n_14747;
or2_13188: n_14740 <=  n_14741  OR n_14744;
and2_13189: n_14741 <=  n_14742  AND n_14743;
inv_13190: n_14742  <= TRANSPORT NOT a_N2348  ;
delay_13191: n_14743  <= TRANSPORT a_SCH3ADDRREG_F3_G  ;
and2_13192: n_14744 <=  n_14745  AND n_14746;
inv_13193: n_14745  <= TRANSPORT NOT a_N2351  ;
delay_13194: n_14746  <= TRANSPORT a_SCH1WRDCNTREG_F3_G  ;
and1_13195: n_14747 <=  gnd;
delay_13196: a_LC2_C8  <= TRANSPORT a_EQ064  ;
xor2_13197: a_EQ064 <=  n_14750  XOR n_14757;
or2_13198: n_14750 <=  n_14751  OR n_14754;
and2_13199: n_14751 <=  n_14752  AND n_14753;
inv_13200: n_14752  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13201: n_14753  <= TRANSPORT a_SCH2ADDRREG_F3_G  ;
and2_13202: n_14754 <=  n_14755  AND n_14756;
inv_13203: n_14755  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13204: n_14756  <= TRANSPORT a_SCH2WRDCNTREG_F3_G  ;
and1_13205: n_14757 <=  gnd;
delay_13206: a_LC1_C8  <= TRANSPORT a_EQ065  ;
xor2_13207: a_EQ065 <=  n_14760  XOR n_14767;
or3_13208: n_14760 <=  n_14761  OR n_14763  OR n_14765;
and1_13209: n_14761 <=  n_14762;
delay_13210: n_14762  <= TRANSPORT a_LC6_C13  ;
and1_13211: n_14763 <=  n_14764;
delay_13212: n_14764  <= TRANSPORT a_LC3_C8  ;
and1_13213: n_14765 <=  n_14766;
delay_13214: n_14766  <= TRANSPORT a_LC2_C8  ;
and1_13215: n_14767 <=  gnd;
delay_13216: a_LC8_C19  <= TRANSPORT a_EQ061  ;
xor2_13217: a_EQ061 <=  n_14770  XOR n_14777;
or2_13218: n_14770 <=  n_14771  OR n_14774;
and2_13219: n_14771 <=  n_14772  AND n_14773;
delay_13220: n_14772  <= TRANSPORT a_N2354_aNOT  ;
delay_13221: n_14773  <= TRANSPORT a_SCH0ADDRREG_F3_G  ;
and2_13222: n_14774 <=  n_14775  AND n_14776;
inv_13223: n_14775  <= TRANSPORT NOT a_N2347  ;
delay_13224: n_14776  <= TRANSPORT a_SCH3WRDCNTREG_F3_G  ;
and1_13225: n_14777 <=  gnd;
delay_13226: a_LC2_A10  <= TRANSPORT a_EQ071  ;
xor2_13227: a_EQ071 <=  n_14780  XOR n_14790;
or3_13228: n_14780 <=  n_14781  OR n_14784  OR n_14787;
and2_13229: n_14781 <=  n_14782  AND n_14783;
delay_13230: n_14782  <= TRANSPORT bytepointer  ;
delay_13231: n_14783  <= TRANSPORT a_LC1_A10  ;
and2_13232: n_14784 <=  n_14785  AND n_14786;
inv_13233: n_14785  <= TRANSPORT NOT bytepointer  ;
delay_13234: n_14786  <= TRANSPORT a_LC1_C8  ;
and2_13235: n_14787 <=  n_14788  AND n_14789;
inv_13236: n_14788  <= TRANSPORT NOT bytepointer  ;
delay_13237: n_14789  <= TRANSPORT a_LC8_C19  ;
and1_13238: n_14790 <=  gnd;
delay_13239: a_LC1_A27  <= TRANSPORT a_EQ072  ;
xor2_13240: a_EQ072 <=  n_14793  XOR n_14799;
or2_13241: n_14793 <=  n_14794  OR n_14796;
and1_13242: n_14794 <=  n_14795;
delay_13243: n_14795  <= TRANSPORT a_LC2_A10  ;
and2_13244: n_14796 <=  n_14797  AND n_14798;
inv_13245: n_14797  <= TRANSPORT NOT a_LC4_A3  ;
delay_13246: n_14798  <= TRANSPORT a_STEMPORARYREG_F3_G  ;
and1_13247: n_14799 <=  gnd;
delay_13248: a_LC5_E10  <= TRANSPORT a_EQ484  ;
xor2_13249: a_EQ484 <=  n_14802  XOR n_14811;
or2_13250: n_14802 <=  n_14803  OR n_14807;
and3_13251: n_14803 <=  n_14804  AND n_14805  AND n_14806;
delay_13252: n_14804  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_13253: n_14805  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_13254: n_14806  <= TRANSPORT a_SCH2MODEREG_F1_G  ;
and3_13255: n_14807 <=  n_14808  AND n_14809  AND n_14810;
inv_13256: n_14808  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_13257: n_14809  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
delay_13258: n_14810  <= TRANSPORT a_SCH1MODEREG_F1_G  ;
and1_13259: n_14811 <=  gnd;
delay_13260: a_LC7_E10  <= TRANSPORT a_EQ485  ;
xor2_13261: a_EQ485 <=  n_14814  XOR n_14823;
or2_13262: n_14814 <=  n_14815  OR n_14819;
and3_13263: n_14815 <=  n_14816  AND n_14817  AND n_14818;
inv_13264: n_14816  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
inv_13265: n_14817  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_13266: n_14818  <= TRANSPORT a_SCH0MODEREG_F1_G  ;
and3_13267: n_14819 <=  n_14820  AND n_14821  AND n_14822;
delay_13268: n_14820  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
delay_13269: n_14821  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
delay_13270: n_14822  <= TRANSPORT a_SCH3MODEREG_F1_G  ;
and1_13271: n_14823 <=  gnd;
delay_13272: a_N1671_aNOT  <= TRANSPORT a_EQ483  ;
xor2_13273: a_EQ483 <=  n_14826  XOR n_14833;
or2_13274: n_14826 <=  n_14827  OR n_14830;
and2_13275: n_14827 <=  n_14828  AND n_14829;
delay_13276: n_14828  <= TRANSPORT a_N66  ;
delay_13277: n_14829  <= TRANSPORT a_LC5_E10  ;
and2_13278: n_14830 <=  n_14831  AND n_14832;
delay_13279: n_14831  <= TRANSPORT a_N66  ;
delay_13280: n_14832  <= TRANSPORT a_LC7_E10  ;
and1_13281: n_14833 <=  gnd;
delay_13282: a_LC4_B7  <= TRANSPORT a_EQ073  ;
xor2_13283: a_EQ073 <=  n_14836  XOR n_14843;
or2_13284: n_14836 <=  n_14837  OR n_14840;
and2_13285: n_14837 <=  n_14838  AND n_14839;
inv_13286: n_14838  <= TRANSPORT NOT a_SMASKREG_F3_G_aNOT  ;
delay_13287: n_14839  <= TRANSPORT a_N2389  ;
and2_13288: n_14840 <=  n_14841  AND n_14842;
inv_13289: n_14841  <= TRANSPORT NOT a_N2367  ;
delay_13290: n_14842  <= TRANSPORT a_STCSTATUS_F3_G  ;
and1_13291: n_14843 <=  gnd;
delay_13292: a_LC2_B18  <= TRANSPORT a_EQ074  ;
xor2_13293: a_EQ074 <=  n_14846  XOR n_14853;
or2_13294: n_14846 <=  n_14847  OR n_14850;
and2_13295: n_14847 <=  n_14848  AND n_14849;
inv_13296: n_14848  <= TRANSPORT NOT a_N63_aNOT  ;
delay_13297: n_14849  <= TRANSPORT a_SREQUESTREG_F3_G  ;
and2_13298: n_14850 <=  n_14851  AND n_14852;
delay_13299: n_14851  <= TRANSPORT a_N73  ;
delay_13300: n_14852  <= TRANSPORT a_SCOMMANDREG_F3_G  ;
and1_13301: n_14853 <=  gnd;
delay_13302: a_LC6_B18  <= TRANSPORT a_EQ075  ;
xor2_13303: a_EQ075 <=  n_14856  XOR n_14863;
or3_13304: n_14856 <=  n_14857  OR n_14859  OR n_14861;
and1_13305: n_14857 <=  n_14858;
delay_13306: n_14858  <= TRANSPORT a_N1671_aNOT  ;
and1_13307: n_14859 <=  n_14860;
delay_13308: n_14860  <= TRANSPORT a_LC4_B7  ;
and1_13309: n_14861 <=  n_14862;
delay_13310: n_14862  <= TRANSPORT a_LC2_B18  ;
and1_13311: n_14863 <=  gnd;
delay_13312: a_G186  <= TRANSPORT a_EQ076  ;
xor2_13313: a_EQ076 <=  n_14865  XOR n_14875;
or3_13314: n_14865 <=  n_14866  OR n_14869  OR n_14872;
and2_13315: n_14866 <=  n_14867  AND n_14868;
inv_13316: n_14867  <= TRANSPORT NOT a_SAEN_aNOT  ;
delay_13317: n_14868  <= TRANSPORT a_LC2_A27  ;
and2_13318: n_14869 <=  n_14870  AND n_14871;
delay_13319: n_14870  <= TRANSPORT a_SAEN_aNOT  ;
delay_13320: n_14871  <= TRANSPORT a_LC1_A27  ;
and2_13321: n_14872 <=  n_14873  AND n_14874;
delay_13322: n_14873  <= TRANSPORT a_SAEN_aNOT  ;
delay_13323: n_14874  <= TRANSPORT a_LC6_B18  ;
and1_13324: n_14875 <=  gnd;
delay_13325: a_LC8_A27  <= TRANSPORT a_EQ139  ;
xor2_13326: a_EQ139 <=  n_14878  XOR n_14887;
or3_13327: n_14878 <=  n_14879  OR n_14882  OR n_14885;
and2_13328: n_14879 <=  n_14880  AND n_14881;
delay_13329: n_14880  <= TRANSPORT a_N1584  ;
delay_13330: n_14881  <= TRANSPORT a_STEMPORARYREG_F4_G  ;
and2_13331: n_14882 <=  n_14883  AND n_14884;
inv_13332: n_14883  <= TRANSPORT NOT a_N1584  ;
delay_13333: n_14884  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and1_13334: n_14885 <=  n_14886;
delay_13335: n_14886  <= TRANSPORT a_SAEN_aNOT  ;
and1_13336: n_14887 <=  gnd;
delay_13337: a_LC5_B7  <= TRANSPORT a_EQ389  ;
xor2_13338: a_EQ389 <=  n_14890  XOR n_14897;
or3_13339: n_14890 <=  n_14891  OR n_14893  OR n_14895;
and1_13340: n_14891 <=  n_14892;
delay_13341: n_14892  <= TRANSPORT a_N2389  ;
and1_13342: n_14893 <=  n_14894;
inv_13343: n_14894  <= TRANSPORT NOT a_N63_aNOT  ;
and1_13344: n_14895 <=  n_14896;
inv_13345: n_14896  <= TRANSPORT NOT a_SAEN_aNOT  ;
and1_13346: n_14897 <=  gnd;
delay_13347: a_LC6_B27  <= TRANSPORT a_EQ486  ;
xor2_13348: a_EQ486 <=  n_14900  XOR n_14909;
or2_13349: n_14900 <=  n_14901  OR n_14905;
and3_13350: n_14901 <=  n_14902  AND n_14903  AND n_14904;
inv_13351: n_14902  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_13352: n_14903  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
delay_13353: n_14904  <= TRANSPORT a_SCH1MODEREG_F2_G  ;
and3_13354: n_14905 <=  n_14906  AND n_14907  AND n_14908;
inv_13355: n_14906  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
inv_13356: n_14907  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_13357: n_14908  <= TRANSPORT a_SCH0MODEREG_F2_G  ;
and1_13358: n_14909 <=  gnd;
delay_13359: a_LC5_B27  <= TRANSPORT a_EQ487  ;
xor2_13360: a_EQ487 <=  n_14912  XOR n_14921;
or2_13361: n_14912 <=  n_14913  OR n_14917;
and3_13362: n_14913 <=  n_14914  AND n_14915  AND n_14916;
delay_13363: n_14914  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
delay_13364: n_14915  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
delay_13365: n_14916  <= TRANSPORT a_SCH3MODEREG_F2_G  ;
and3_13366: n_14917 <=  n_14918  AND n_14919  AND n_14920;
delay_13367: n_14918  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_13368: n_14919  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_13369: n_14920  <= TRANSPORT a_SCH2MODEREG_F2_G  ;
and1_13370: n_14921 <=  gnd;
delay_13371: a_N1693_aNOT  <= TRANSPORT a_EQ488  ;
xor2_13372: a_EQ488 <=  n_14924  XOR n_14931;
or2_13373: n_14924 <=  n_14925  OR n_14928;
and2_13374: n_14925 <=  n_14926  AND n_14927;
delay_13375: n_14926  <= TRANSPORT a_N66  ;
delay_13376: n_14927  <= TRANSPORT a_LC6_B27  ;
and2_13377: n_14928 <=  n_14929  AND n_14930;
delay_13378: n_14929  <= TRANSPORT a_N66  ;
delay_13379: n_14930  <= TRANSPORT a_LC5_B27  ;
and1_13380: n_14931 <=  gnd;
delay_13381: a_LC1_B27  <= TRANSPORT a_EQ140  ;
xor2_13382: a_EQ140 <=  n_14934  XOR n_14940;
or2_13383: n_14934 <=  n_14935  OR n_14937;
and1_13384: n_14935 <=  n_14936;
delay_13385: n_14936  <= TRANSPORT a_N1693_aNOT  ;
and2_13386: n_14937 <=  n_14938  AND n_14939;
delay_13387: n_14938  <= TRANSPORT a_N73  ;
delay_13388: n_14939  <= TRANSPORT a_SCOMMANDREG_F4_G  ;
and1_13389: n_14940 <=  gnd;
delay_13390: a_LC8_B14  <= TRANSPORT a_EQ137  ;
xor2_13391: a_EQ137 <=  n_14943  XOR n_14952;
or2_13392: n_14943 <=  n_14944  OR n_14948;
and3_13393: n_14944 <=  n_14945  AND n_14946  AND n_14947;
inv_13394: n_14945  <= TRANSPORT NOT a_N2367  ;
delay_13395: n_14946  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
inv_13396: n_14947  <= TRANSPORT NOT a_N4185  ;
and3_13397: n_14948 <=  n_14949  AND n_14950  AND n_14951;
inv_13398: n_14949  <= TRANSPORT NOT a_N2367  ;
inv_13399: n_14950  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
delay_13400: n_14951  <= TRANSPORT a_N4185  ;
and1_13401: n_14952 <=  gnd;
delay_13402: a_LC1_C19  <= TRANSPORT a_EQ127  ;
xor2_13403: a_EQ127 <=  n_14955  XOR n_14962;
or2_13404: n_14955 <=  n_14956  OR n_14959;
and2_13405: n_14956 <=  n_14957  AND n_14958;
inv_13406: n_14957  <= TRANSPORT NOT a_N2353  ;
delay_13407: n_14958  <= TRANSPORT a_SCH0WRDCNTREG_F4_G  ;
and2_13408: n_14959 <=  n_14960  AND n_14961;
inv_13409: n_14960  <= TRANSPORT NOT a_N2347  ;
delay_13410: n_14961  <= TRANSPORT a_SCH3WRDCNTREG_F4_G  ;
and1_13411: n_14962 <=  gnd;
delay_13412: a_LC4_C19  <= TRANSPORT a_EQ128  ;
xor2_13413: a_EQ128 <=  n_14965  XOR n_14972;
or2_13414: n_14965 <=  n_14966  OR n_14969;
and2_13415: n_14966 <=  n_14967  AND n_14968;
inv_13416: n_14967  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13417: n_14968  <= TRANSPORT a_SCH2ADDRREG_F4_G  ;
and2_13418: n_14969 <=  n_14970  AND n_14971;
inv_13419: n_14970  <= TRANSPORT NOT a_N2352  ;
delay_13420: n_14971  <= TRANSPORT a_SCH1ADDRREG_F4_G  ;
and1_13421: n_14972 <=  gnd;
delay_13422: a_LC5_C19  <= TRANSPORT a_EQ129  ;
xor2_13423: a_EQ129 <=  n_14975  XOR n_14982;
or2_13424: n_14975 <=  n_14976  OR n_14979;
and2_13425: n_14976 <=  n_14977  AND n_14978;
inv_13426: n_14977  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13427: n_14978  <= TRANSPORT a_SCH2WRDCNTREG_F4_G  ;
and2_13428: n_14979 <=  n_14980  AND n_14981;
inv_13429: n_14980  <= TRANSPORT NOT a_N2348  ;
delay_13430: n_14981  <= TRANSPORT a_SCH3ADDRREG_F4_G  ;
and1_13431: n_14982 <=  gnd;
delay_13432: a_LC6_C19  <= TRANSPORT a_EQ130  ;
xor2_13433: a_EQ130 <=  n_14985  XOR n_14992;
or2_13434: n_14985 <=  n_14986  OR n_14989;
and2_13435: n_14986 <=  n_14987  AND n_14988;
delay_13436: n_14987  <= TRANSPORT a_N2354_aNOT  ;
delay_13437: n_14988  <= TRANSPORT a_SCH0ADDRREG_F4_G  ;
and2_13438: n_14989 <=  n_14990  AND n_14991;
inv_13439: n_14990  <= TRANSPORT NOT a_N2351  ;
delay_13440: n_14991  <= TRANSPORT a_SCH1WRDCNTREG_F4_G  ;
and1_13441: n_14992 <=  gnd;
delay_13442: a_LC2_C19  <= TRANSPORT a_EQ131  ;
xor2_13443: a_EQ131 <=  n_14995  XOR n_15004;
or4_13444: n_14995 <=  n_14996  OR n_14998  OR n_15000  OR n_15002;
and1_13445: n_14996 <=  n_14997;
delay_13446: n_14997  <= TRANSPORT a_LC1_C19  ;
and1_13447: n_14998 <=  n_14999;
delay_13448: n_14999  <= TRANSPORT a_LC4_C19  ;
and1_13449: n_15000 <=  n_15001;
delay_13450: n_15001  <= TRANSPORT a_LC5_C19  ;
and1_13451: n_15002 <=  n_15003;
delay_13452: n_15003  <= TRANSPORT a_LC6_C19  ;
and1_13453: n_15004 <=  gnd;
delay_13454: a_LC6_A6  <= TRANSPORT a_EQ132  ;
xor2_13455: a_EQ132 <=  n_15007  XOR n_15014;
or2_13456: n_15007 <=  n_15008  OR n_15011;
and2_13457: n_15008 <=  n_15009  AND n_15010;
inv_13458: n_15009  <= TRANSPORT NOT a_N2353  ;
delay_13459: n_15010  <= TRANSPORT a_SH0WRDCNTREG_F12_G  ;
and2_13460: n_15011 <=  n_15012  AND n_15013;
inv_13461: n_15012  <= TRANSPORT NOT a_N2347  ;
delay_13462: n_15013  <= TRANSPORT a_SH3WRDCNTREG_F12_G  ;
and1_13463: n_15014 <=  gnd;
delay_13464: a_LC5_A6  <= TRANSPORT a_EQ133  ;
xor2_13465: a_EQ133 <=  n_15017  XOR n_15024;
or2_13466: n_15017 <=  n_15018  OR n_15021;
and2_13467: n_15018 <=  n_15019  AND n_15020;
inv_13468: n_15019  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13469: n_15020  <= TRANSPORT a_SCH2ADDRREG_F12_G  ;
and2_13470: n_15021 <=  n_15022  AND n_15023;
inv_13471: n_15022  <= TRANSPORT NOT a_N2352  ;
delay_13472: n_15023  <= TRANSPORT a_SCH1ADDRREG_F12_G  ;
and1_13473: n_15024 <=  gnd;
delay_13474: a_LC4_A6  <= TRANSPORT a_EQ134  ;
xor2_13475: a_EQ134 <=  n_15027  XOR n_15034;
or2_13476: n_15027 <=  n_15028  OR n_15031;
and2_13477: n_15028 <=  n_15029  AND n_15030;
inv_13478: n_15029  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13479: n_15030  <= TRANSPORT a_SH2WRDCNTREG_F12_G  ;
and2_13480: n_15031 <=  n_15032  AND n_15033;
inv_13481: n_15032  <= TRANSPORT NOT a_N2348  ;
delay_13482: n_15033  <= TRANSPORT a_SCH3ADDRREG_F12_G  ;
and1_13483: n_15034 <=  gnd;
delay_13484: a_LC3_A6  <= TRANSPORT a_EQ135  ;
xor2_13485: a_EQ135 <=  n_15037  XOR n_15044;
or2_13486: n_15037 <=  n_15038  OR n_15041;
and2_13487: n_15038 <=  n_15039  AND n_15040;
delay_13488: n_15039  <= TRANSPORT a_N2354_aNOT  ;
delay_13489: n_15040  <= TRANSPORT a_SCH0ADDRREG_F12_G  ;
and2_13490: n_15041 <=  n_15042  AND n_15043;
inv_13491: n_15042  <= TRANSPORT NOT a_N2351  ;
delay_13492: n_15043  <= TRANSPORT a_SH1WRDCNTREG_F12_G  ;
and1_13493: n_15044 <=  gnd;
delay_13494: a_LC2_A6  <= TRANSPORT a_EQ136  ;
xor2_13495: a_EQ136 <=  n_15047  XOR n_15056;
or4_13496: n_15047 <=  n_15048  OR n_15050  OR n_15052  OR n_15054;
and1_13497: n_15048 <=  n_15049;
delay_13498: n_15049  <= TRANSPORT a_LC6_A6  ;
and1_13499: n_15050 <=  n_15051;
delay_13500: n_15051  <= TRANSPORT a_LC5_A6  ;
and1_13501: n_15052 <=  n_15053;
delay_13502: n_15053  <= TRANSPORT a_LC4_A6  ;
and1_13503: n_15054 <=  n_15055;
delay_13504: n_15055  <= TRANSPORT a_LC3_A6  ;
and1_13505: n_15056 <=  gnd;
delay_13506: a_LC1_A6  <= TRANSPORT a_EQ138  ;
xor2_13507: a_EQ138 <=  n_15059  XOR n_15068;
or3_13508: n_15059 <=  n_15060  OR n_15062  OR n_15065;
and1_13509: n_15060 <=  n_15061;
delay_13510: n_15061  <= TRANSPORT a_LC8_B14  ;
and2_13511: n_15062 <=  n_15063  AND n_15064;
inv_13512: n_15063  <= TRANSPORT NOT bytepointer  ;
delay_13513: n_15064  <= TRANSPORT a_LC2_C19  ;
and2_13514: n_15065 <=  n_15066  AND n_15067;
delay_13515: n_15066  <= TRANSPORT bytepointer  ;
delay_13516: n_15067  <= TRANSPORT a_LC2_A6  ;
and1_13517: n_15068 <=  gnd;
delay_13518: a_LC7_A27  <= TRANSPORT a_EQ141  ;
xor2_13519: a_EQ141 <=  n_15071  XOR n_15081;
or3_13520: n_15071 <=  n_15072  OR n_15075  OR n_15078;
and2_13521: n_15072 <=  n_15073  AND n_15074;
delay_13522: n_15073  <= TRANSPORT a_LC8_A27  ;
delay_13523: n_15074  <= TRANSPORT a_LC5_B7  ;
and2_13524: n_15075 <=  n_15076  AND n_15077;
delay_13525: n_15076  <= TRANSPORT a_LC8_A27  ;
delay_13526: n_15077  <= TRANSPORT a_LC1_B27  ;
and2_13527: n_15078 <=  n_15079  AND n_15080;
delay_13528: n_15079  <= TRANSPORT a_LC8_A27  ;
delay_13529: n_15080  <= TRANSPORT a_LC1_A6  ;
and1_13530: n_15081 <=  gnd;
delay_13531: a_LC6_A27  <= TRANSPORT a_EQ126  ;
xor2_13532: a_EQ126 <=  n_15084  XOR n_15091;
or3_13533: n_15084 <=  n_15085  OR n_15087  OR n_15089;
and1_13534: n_15085 <=  n_15086;
delay_13535: n_15086  <= TRANSPORT a_SAEN_aNOT  ;
and1_13536: n_15087 <=  n_15088;
delay_13537: n_15088  <= TRANSPORT a_SADDRESSOUT_F12_G  ;
and1_13538: n_15089 <=  n_15090;
delay_13539: n_15090  <= TRANSPORT a_N1584  ;
and1_13540: n_15091 <=  gnd;
delay_13541: a_G993  <= TRANSPORT a_EQ142  ;
xor2_13542: a_EQ142 <=  n_15093  XOR n_15100;
or2_13543: n_15093 <=  n_15094  OR n_15096;
and1_13544: n_15094 <=  n_15095;
delay_13545: n_15095  <= TRANSPORT a_LC7_A27  ;
and3_13546: n_15096 <=  n_15097  AND n_15098  AND n_15099;
inv_13547: n_15097  <= TRANSPORT NOT a_LC4_A3  ;
delay_13548: n_15098  <= TRANSPORT a_STEMPORARYREG_F4_G  ;
delay_13549: n_15099  <= TRANSPORT a_LC6_A27  ;
and1_13550: n_15100 <=  gnd;
delay_13551: a_LC6_E1  <= TRANSPORT a_EQ510  ;
xor2_13552: a_EQ510 <=  n_15103  XOR n_15112;
or2_13553: n_15103 <=  n_15104  OR n_15108;
and3_13554: n_15104 <=  n_15105  AND n_15106  AND n_15107;
delay_13555: n_15105  <= TRANSPORT a_SCH2MODEREG_F3_G  ;
delay_13556: n_15106  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_13557: n_15107  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and3_13558: n_15108 <=  n_15109  AND n_15110  AND n_15111;
delay_13559: n_15109  <= TRANSPORT a_SCH0MODEREG_F3_G  ;
inv_13560: n_15110  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
inv_13561: n_15111  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and1_13562: n_15112 <=  gnd;
delay_13563: a_LC5_E1  <= TRANSPORT a_EQ511  ;
xor2_13564: a_EQ511 <=  n_15115  XOR n_15124;
or2_13565: n_15115 <=  n_15116  OR n_15120;
and3_13566: n_15116 <=  n_15117  AND n_15118  AND n_15119;
delay_13567: n_15117  <= TRANSPORT a_SCH1MODEREG_F3_G  ;
inv_13568: n_15118  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_13569: n_15119  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and3_13570: n_15120 <=  n_15121  AND n_15122  AND n_15123;
delay_13571: n_15121  <= TRANSPORT a_SCH3MODEREG_F3_G  ;
delay_13572: n_15122  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
delay_13573: n_15123  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and1_13574: n_15124 <=  gnd;
delay_13575: a_N1837_aNOT  <= TRANSPORT a_EQ509  ;
xor2_13576: a_EQ509 <=  n_15127  XOR n_15134;
or2_13577: n_15127 <=  n_15128  OR n_15131;
and2_13578: n_15128 <=  n_15129  AND n_15130;
delay_13579: n_15129  <= TRANSPORT a_N66  ;
delay_13580: n_15130  <= TRANSPORT a_LC6_E1  ;
and2_13581: n_15131 <=  n_15132  AND n_15133;
delay_13582: n_15132  <= TRANSPORT a_N66  ;
delay_13583: n_15133  <= TRANSPORT a_LC5_E1  ;
and1_13584: n_15134 <=  gnd;
delay_13585: a_LC8_F11  <= TRANSPORT a_EQ095  ;
xor2_13586: a_EQ095 <=  n_15137  XOR n_15144;
or2_13587: n_15137 <=  n_15138  OR n_15141;
and2_13588: n_15138 <=  n_15139  AND n_15140;
inv_13589: n_15139  <= TRANSPORT NOT a_N2353  ;
delay_13590: n_15140  <= TRANSPORT a_SCH0WRDCNTREG_F5_G  ;
and2_13591: n_15141 <=  n_15142  AND n_15143;
inv_13592: n_15142  <= TRANSPORT NOT a_N2347  ;
delay_13593: n_15143  <= TRANSPORT a_SCH3WRDCNTREG_F5_G  ;
and1_13594: n_15144 <=  gnd;
delay_13595: a_LC7_F11  <= TRANSPORT a_EQ096  ;
xor2_13596: a_EQ096 <=  n_15147  XOR n_15154;
or2_13597: n_15147 <=  n_15148  OR n_15151;
and2_13598: n_15148 <=  n_15149  AND n_15150;
inv_13599: n_15149  <= TRANSPORT NOT a_N2351  ;
delay_13600: n_15150  <= TRANSPORT a_SCH1WRDCNTREG_F5_G  ;
and2_13601: n_15151 <=  n_15152  AND n_15153;
inv_13602: n_15152  <= TRANSPORT NOT a_N2352  ;
delay_13603: n_15153  <= TRANSPORT a_SCH1ADDRREG_F5_G  ;
and1_13604: n_15154 <=  gnd;
delay_13605: a_LC6_F19  <= TRANSPORT a_EQ097  ;
xor2_13606: a_EQ097 <=  n_15157  XOR n_15164;
or2_13607: n_15157 <=  n_15158  OR n_15161;
and2_13608: n_15158 <=  n_15159  AND n_15160;
inv_13609: n_15159  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13610: n_15160  <= TRANSPORT a_SCH2WRDCNTREG_F5_G  ;
and2_13611: n_15161 <=  n_15162  AND n_15163;
inv_13612: n_15162  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13613: n_15163  <= TRANSPORT a_SCH2ADDRREG_F5_G  ;
and1_13614: n_15164 <=  gnd;
delay_13615: a_LC6_F11  <= TRANSPORT a_EQ098  ;
xor2_13616: a_EQ098 <=  n_15167  XOR n_15174;
or2_13617: n_15167 <=  n_15168  OR n_15171;
and2_13618: n_15168 <=  n_15169  AND n_15170;
delay_13619: n_15169  <= TRANSPORT a_N2354_aNOT  ;
delay_13620: n_15170  <= TRANSPORT a_SCH0ADDRREG_F5_G  ;
and2_13621: n_15171 <=  n_15172  AND n_15173;
inv_13622: n_15172  <= TRANSPORT NOT a_N2348  ;
delay_13623: n_15173  <= TRANSPORT a_SCH3ADDRREG_F5_G  ;
and1_13624: n_15174 <=  gnd;
delay_13625: a_LC3_F11  <= TRANSPORT a_EQ099  ;
xor2_13626: a_EQ099 <=  n_15177  XOR n_15186;
or4_13627: n_15177 <=  n_15178  OR n_15180  OR n_15182  OR n_15184;
and1_13628: n_15178 <=  n_15179;
delay_13629: n_15179  <= TRANSPORT a_LC8_F11  ;
and1_13630: n_15180 <=  n_15181;
delay_13631: n_15181  <= TRANSPORT a_LC7_F11  ;
and1_13632: n_15182 <=  n_15183;
delay_13633: n_15183  <= TRANSPORT a_LC6_F19  ;
and1_13634: n_15184 <=  n_15185;
delay_13635: n_15185  <= TRANSPORT a_LC6_F11  ;
and1_13636: n_15186 <=  gnd;
delay_13637: a_LC7_E7  <= TRANSPORT a_EQ100  ;
xor2_13638: a_EQ100 <=  n_15189  XOR n_15196;
or2_13639: n_15189 <=  n_15190  OR n_15193;
and2_13640: n_15190 <=  n_15191  AND n_15192;
inv_13641: n_15191  <= TRANSPORT NOT a_N2353  ;
delay_13642: n_15192  <= TRANSPORT a_SH0WRDCNTREG_F13_G  ;
and2_13643: n_15193 <=  n_15194  AND n_15195;
inv_13644: n_15194  <= TRANSPORT NOT a_N2347  ;
delay_13645: n_15195  <= TRANSPORT a_SH3WRDCNTREG_F13_G  ;
and1_13646: n_15196 <=  gnd;
delay_13647: a_LC6_E7  <= TRANSPORT a_EQ101  ;
xor2_13648: a_EQ101 <=  n_15199  XOR n_15206;
or2_13649: n_15199 <=  n_15200  OR n_15203;
and2_13650: n_15200 <=  n_15201  AND n_15202;
inv_13651: n_15201  <= TRANSPORT NOT a_N2351  ;
delay_13652: n_15202  <= TRANSPORT a_SH1WRDCNTREG_F13_G  ;
and2_13653: n_15203 <=  n_15204  AND n_15205;
inv_13654: n_15204  <= TRANSPORT NOT a_N2352  ;
delay_13655: n_15205  <= TRANSPORT a_SCH1ADDRREG_F13_G  ;
and1_13656: n_15206 <=  gnd;
delay_13657: a_LC5_E7  <= TRANSPORT a_EQ102  ;
xor2_13658: a_EQ102 <=  n_15209  XOR n_15216;
or2_13659: n_15209 <=  n_15210  OR n_15213;
and2_13660: n_15210 <=  n_15211  AND n_15212;
inv_13661: n_15211  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13662: n_15212  <= TRANSPORT a_SH2WRDCNTREG_F13_G  ;
and2_13663: n_15213 <=  n_15214  AND n_15215;
inv_13664: n_15214  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13665: n_15215  <= TRANSPORT a_SCH2ADDRREG_F13_G  ;
and1_13666: n_15216 <=  gnd;
delay_13667: a_LC2_E14  <= TRANSPORT a_EQ103  ;
xor2_13668: a_EQ103 <=  n_15219  XOR n_15226;
or2_13669: n_15219 <=  n_15220  OR n_15223;
and2_13670: n_15220 <=  n_15221  AND n_15222;
delay_13671: n_15221  <= TRANSPORT a_N2354_aNOT  ;
delay_13672: n_15222  <= TRANSPORT a_SCH0ADDRREG_F13_G  ;
and2_13673: n_15223 <=  n_15224  AND n_15225;
inv_13674: n_15224  <= TRANSPORT NOT a_N2348  ;
delay_13675: n_15225  <= TRANSPORT a_SCH3ADDRREG_F13_G  ;
and1_13676: n_15226 <=  gnd;
delay_13677: a_LC4_E7  <= TRANSPORT a_EQ104  ;
xor2_13678: a_EQ104 <=  n_15229  XOR n_15238;
or4_13679: n_15229 <=  n_15230  OR n_15232  OR n_15234  OR n_15236;
and1_13680: n_15230 <=  n_15231;
delay_13681: n_15231  <= TRANSPORT a_LC7_E7  ;
and1_13682: n_15232 <=  n_15233;
delay_13683: n_15233  <= TRANSPORT a_LC6_E7  ;
and1_13684: n_15234 <=  n_15235;
delay_13685: n_15235  <= TRANSPORT a_LC5_E7  ;
and1_13686: n_15236 <=  n_15237;
delay_13687: n_15237  <= TRANSPORT a_LC2_E14  ;
and1_13688: n_15238 <=  gnd;
delay_13689: a_LC3_E7  <= TRANSPORT a_EQ105  ;
xor2_13690: a_EQ105 <=  n_15241  XOR n_15250;
or3_13691: n_15241 <=  n_15242  OR n_15244  OR n_15247;
and1_13692: n_15242 <=  n_15243;
delay_13693: n_15243  <= TRANSPORT a_N1837_aNOT  ;
and2_13694: n_15244 <=  n_15245  AND n_15246;
inv_13695: n_15245  <= TRANSPORT NOT bytepointer  ;
delay_13696: n_15246  <= TRANSPORT a_LC3_F11  ;
and2_13697: n_15247 <=  n_15248  AND n_15249;
delay_13698: n_15248  <= TRANSPORT bytepointer  ;
delay_13699: n_15249  <= TRANSPORT a_LC4_E7  ;
and1_13700: n_15250 <=  gnd;
delay_13701: a_N1849  <= TRANSPORT a_N1849_aIN  ;
xor2_13702: a_N1849_aIN <=  n_15253  XOR n_15257;
or1_13703: n_15253 <=  n_15254;
and2_13704: n_15254 <=  n_15255  AND n_15256;
inv_13705: n_15255  <= TRANSPORT NOT a_N2557  ;
delay_13706: n_15256  <= TRANSPORT a_SADDRESSOUT_F13_G  ;
and1_13707: n_15257 <=  gnd;
delay_13708: a_LC2_E7  <= TRANSPORT a_EQ106  ;
xor2_13709: a_EQ106 <=  n_15260  XOR n_15268;
or3_13710: n_15260 <=  n_15261  OR n_15263  OR n_15266;
and1_13711: n_15261 <=  n_15262;
delay_13712: n_15262  <= TRANSPORT a_N1849  ;
and2_13713: n_15263 <=  n_15264  AND n_15265;
delay_13714: n_15264  <= TRANSPORT a_N1584  ;
delay_13715: n_15265  <= TRANSPORT a_STEMPORARYREG_F5_G  ;
and1_13716: n_15266 <=  n_15267;
delay_13717: n_15267  <= TRANSPORT a_SAEN_aNOT  ;
and1_13718: n_15268 <=  gnd;
delay_13719: a_LC6_B24  <= TRANSPORT a_EQ107  ;
xor2_13720: a_EQ107 <=  n_15271  XOR n_15278;
or2_13721: n_15271 <=  n_15272  OR n_15275;
and2_13722: n_15272 <=  n_15273  AND n_15274;
delay_13723: n_15273  <= TRANSPORT a_STEMPORARYREG_F5_G  ;
delay_13724: n_15274  <= TRANSPORT a_N1830  ;
and2_13725: n_15275 <=  n_15276  AND n_15277;
delay_13726: n_15276  <= TRANSPORT a_N73  ;
delay_13727: n_15277  <= TRANSPORT a_SCOMMANDREG_F5_G  ;
and1_13728: n_15278 <=  gnd;
delay_13729: a_LC2_B24  <= TRANSPORT a_EQ108  ;
xor2_13730: a_EQ108 <=  n_15281  XOR n_15292;
or3_13731: n_15281 <=  n_15282  OR n_15284  OR n_15288;
and1_13732: n_15282 <=  n_15283;
delay_13733: n_15283  <= TRANSPORT a_LC6_B24  ;
and3_13734: n_15284 <=  n_15285  AND n_15286  AND n_15287;
inv_13735: n_15285  <= TRANSPORT NOT a_N2367  ;
delay_13736: n_15286  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
inv_13737: n_15287  <= TRANSPORT NOT a_N4184  ;
and3_13738: n_15288 <=  n_15289  AND n_15290  AND n_15291;
inv_13739: n_15289  <= TRANSPORT NOT a_N2367  ;
inv_13740: n_15290  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
delay_13741: n_15291  <= TRANSPORT a_N4184  ;
and1_13742: n_15292 <=  gnd;
delay_13743: a_G917  <= TRANSPORT a_EQ109  ;
xor2_13744: a_EQ109 <=  n_15294  XOR n_15304;
or3_13745: n_15294 <=  n_15295  OR n_15298  OR n_15301;
and2_13746: n_15295 <=  n_15296  AND n_15297;
delay_13747: n_15296  <= TRANSPORT a_LC3_E7  ;
delay_13748: n_15297  <= TRANSPORT a_LC2_E7  ;
and2_13749: n_15298 <=  n_15299  AND n_15300;
delay_13750: n_15299  <= TRANSPORT a_LC2_E7  ;
delay_13751: n_15300  <= TRANSPORT a_LC2_B24  ;
and2_13752: n_15301 <=  n_15302  AND n_15303;
delay_13753: n_15302  <= TRANSPORT a_LC5_B7  ;
delay_13754: n_15303  <= TRANSPORT a_LC2_E7  ;
and1_13755: n_15304 <=  gnd;
delay_13756: a_LC5_B14  <= TRANSPORT a_EQ055  ;
xor2_13757: a_EQ055 <=  n_15307  XOR n_15319;
or3_13758: n_15307 <=  n_15308  OR n_15312  OR n_15316;
and3_13759: n_15308 <=  n_15309  AND n_15310  AND n_15311;
inv_13760: n_15309  <= TRANSPORT NOT a_N2367  ;
inv_13761: n_15310  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
delay_13762: n_15311  <= TRANSPORT a_N4183  ;
and3_13763: n_15312 <=  n_15313  AND n_15314  AND n_15315;
inv_13764: n_15313  <= TRANSPORT NOT a_N2367  ;
delay_13765: n_15314  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
inv_13766: n_15315  <= TRANSPORT NOT a_N4183  ;
and2_13767: n_15316 <=  n_15317  AND n_15318;
delay_13768: n_15317  <= TRANSPORT a_N73  ;
delay_13769: n_15318  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
and1_13770: n_15319 <=  gnd;
delay_13771: a_LC7_E18  <= TRANSPORT a_EQ045  ;
xor2_13772: a_EQ045 <=  n_15322  XOR n_15329;
or2_13773: n_15322 <=  n_15323  OR n_15326;
and2_13774: n_15323 <=  n_15324  AND n_15325;
inv_13775: n_15324  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13776: n_15325  <= TRANSPORT a_SH2WRDCNTREG_F14_G  ;
and2_13777: n_15326 <=  n_15327  AND n_15328;
inv_13778: n_15327  <= TRANSPORT NOT a_N2347  ;
delay_13779: n_15328  <= TRANSPORT a_SH3WRDCNTREG_F14_G  ;
and1_13780: n_15329 <=  gnd;
delay_13781: a_LC7_F19  <= TRANSPORT a_EQ046  ;
xor2_13782: a_EQ046 <=  n_15332  XOR n_15339;
or2_13783: n_15332 <=  n_15333  OR n_15336;
and2_13784: n_15333 <=  n_15334  AND n_15335;
inv_13785: n_15334  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13786: n_15335  <= TRANSPORT a_SCH2ADDRREG_F14_G  ;
and2_13787: n_15336 <=  n_15337  AND n_15338;
inv_13788: n_15337  <= TRANSPORT NOT a_N2348  ;
delay_13789: n_15338  <= TRANSPORT a_SCH3ADDRREG_F14_G  ;
and1_13790: n_15339 <=  gnd;
delay_13791: a_LC6_E18  <= TRANSPORT a_EQ047  ;
xor2_13792: a_EQ047 <=  n_15342  XOR n_15349;
or2_13793: n_15342 <=  n_15343  OR n_15346;
and2_13794: n_15343 <=  n_15344  AND n_15345;
inv_13795: n_15344  <= TRANSPORT NOT a_N2351  ;
delay_13796: n_15345  <= TRANSPORT a_SH1WRDCNTREG_F14_G  ;
and2_13797: n_15346 <=  n_15347  AND n_15348;
delay_13798: n_15347  <= TRANSPORT a_N2354_aNOT  ;
delay_13799: n_15348  <= TRANSPORT a_SCH0ADDRREG_F14_G  ;
and1_13800: n_15349 <=  gnd;
delay_13801: a_LC5_E18  <= TRANSPORT a_EQ048  ;
xor2_13802: a_EQ048 <=  n_15352  XOR n_15359;
or2_13803: n_15352 <=  n_15353  OR n_15356;
and2_13804: n_15353 <=  n_15354  AND n_15355;
inv_13805: n_15354  <= TRANSPORT NOT a_N2352  ;
delay_13806: n_15355  <= TRANSPORT a_SCH1ADDRREG_F14_G  ;
and2_13807: n_15356 <=  n_15357  AND n_15358;
inv_13808: n_15357  <= TRANSPORT NOT a_N2353  ;
delay_13809: n_15358  <= TRANSPORT a_SH0WRDCNTREG_F14_G  ;
and1_13810: n_15359 <=  gnd;
delay_13811: a_LC4_E18  <= TRANSPORT a_EQ049  ;
xor2_13812: a_EQ049 <=  n_15362  XOR n_15371;
or4_13813: n_15362 <=  n_15363  OR n_15365  OR n_15367  OR n_15369;
and1_13814: n_15363 <=  n_15364;
delay_13815: n_15364  <= TRANSPORT a_LC7_E18  ;
and1_13816: n_15365 <=  n_15366;
delay_13817: n_15366  <= TRANSPORT a_LC7_F19  ;
and1_13818: n_15367 <=  n_15368;
delay_13819: n_15368  <= TRANSPORT a_LC6_E18  ;
and1_13820: n_15369 <=  n_15370;
delay_13821: n_15370  <= TRANSPORT a_LC5_E18  ;
and1_13822: n_15371 <=  gnd;
delay_13823: a_LC5_F11  <= TRANSPORT a_EQ050  ;
xor2_13824: a_EQ050 <=  n_15374  XOR n_15381;
or2_13825: n_15374 <=  n_15375  OR n_15378;
and2_13826: n_15375 <=  n_15376  AND n_15377;
inv_13827: n_15376  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13828: n_15377  <= TRANSPORT a_SCH2WRDCNTREG_F6_G  ;
and2_13829: n_15378 <=  n_15379  AND n_15380;
inv_13830: n_15379  <= TRANSPORT NOT a_N2347  ;
delay_13831: n_15380  <= TRANSPORT a_SCH3WRDCNTREG_F6_G  ;
and1_13832: n_15381 <=  gnd;
delay_13833: a_LC3_F26  <= TRANSPORT a_EQ051  ;
xor2_13834: a_EQ051 <=  n_15384  XOR n_15391;
or2_13835: n_15384 <=  n_15385  OR n_15388;
and2_13836: n_15385 <=  n_15386  AND n_15387;
inv_13837: n_15386  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13838: n_15387  <= TRANSPORT a_SCH2ADDRREG_F6_G  ;
and2_13839: n_15388 <=  n_15389  AND n_15390;
inv_13840: n_15389  <= TRANSPORT NOT a_N2348  ;
delay_13841: n_15390  <= TRANSPORT a_SCH3ADDRREG_F6_G  ;
and1_13842: n_15391 <=  gnd;
delay_13843: a_LC4_F11  <= TRANSPORT a_EQ052  ;
xor2_13844: a_EQ052 <=  n_15394  XOR n_15401;
or2_13845: n_15394 <=  n_15395  OR n_15398;
and2_13846: n_15395 <=  n_15396  AND n_15397;
inv_13847: n_15396  <= TRANSPORT NOT a_N2351  ;
delay_13848: n_15397  <= TRANSPORT a_SCH1WRDCNTREG_F6_G  ;
and2_13849: n_15398 <=  n_15399  AND n_15400;
delay_13850: n_15399  <= TRANSPORT a_N2354_aNOT  ;
delay_13851: n_15400  <= TRANSPORT a_SCH0ADDRREG_F6_G  ;
and1_13852: n_15401 <=  gnd;
delay_13853: a_LC2_F11  <= TRANSPORT a_EQ053  ;
xor2_13854: a_EQ053 <=  n_15404  XOR n_15411;
or2_13855: n_15404 <=  n_15405  OR n_15408;
and2_13856: n_15405 <=  n_15406  AND n_15407;
inv_13857: n_15406  <= TRANSPORT NOT a_N2352  ;
delay_13858: n_15407  <= TRANSPORT a_SCH1ADDRREG_F6_G  ;
and2_13859: n_15408 <=  n_15409  AND n_15410;
inv_13860: n_15409  <= TRANSPORT NOT a_N2353  ;
delay_13861: n_15410  <= TRANSPORT a_SCH0WRDCNTREG_F6_G  ;
and1_13862: n_15411 <=  gnd;
delay_13863: a_LC1_F11  <= TRANSPORT a_EQ054  ;
xor2_13864: a_EQ054 <=  n_15414  XOR n_15423;
or4_13865: n_15414 <=  n_15415  OR n_15417  OR n_15419  OR n_15421;
and1_13866: n_15415 <=  n_15416;
delay_13867: n_15416  <= TRANSPORT a_LC5_F11  ;
and1_13868: n_15417 <=  n_15418;
delay_13869: n_15418  <= TRANSPORT a_LC3_F26  ;
and1_13870: n_15419 <=  n_15420;
delay_13871: n_15420  <= TRANSPORT a_LC4_F11  ;
and1_13872: n_15421 <=  n_15422;
delay_13873: n_15422  <= TRANSPORT a_LC2_F11  ;
and1_13874: n_15423 <=  gnd;
delay_13875: a_LC3_E18  <= TRANSPORT a_EQ056  ;
xor2_13876: a_EQ056 <=  n_15426  XOR n_15435;
or3_13877: n_15426 <=  n_15427  OR n_15429  OR n_15432;
and1_13878: n_15427 <=  n_15428;
delay_13879: n_15428  <= TRANSPORT a_LC5_B14  ;
and2_13880: n_15429 <=  n_15430  AND n_15431;
delay_13881: n_15430  <= TRANSPORT bytepointer  ;
delay_13882: n_15431  <= TRANSPORT a_LC4_E18  ;
and2_13883: n_15432 <=  n_15433  AND n_15434;
inv_13884: n_15433  <= TRANSPORT NOT bytepointer  ;
delay_13885: n_15434  <= TRANSPORT a_LC1_F11  ;
and1_13886: n_15435 <=  gnd;
delay_13887: a_LC8_E2  <= TRANSPORT a_EQ499  ;
xor2_13888: a_EQ499 <=  n_15438  XOR n_15447;
or2_13889: n_15438 <=  n_15439  OR n_15443;
and3_13890: n_15439 <=  n_15440  AND n_15441  AND n_15442;
delay_13891: n_15440  <= TRANSPORT a_SCH1MODEREG_F4_G  ;
inv_13892: n_15441  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_13893: n_15442  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and3_13894: n_15443 <=  n_15444  AND n_15445  AND n_15446;
delay_13895: n_15444  <= TRANSPORT a_SCH2MODEREG_F4_G  ;
delay_13896: n_15445  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_13897: n_15446  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and1_13898: n_15447 <=  gnd;
delay_13899: a_LC7_E2  <= TRANSPORT a_EQ500  ;
xor2_13900: a_EQ500 <=  n_15450  XOR n_15459;
or2_13901: n_15450 <=  n_15451  OR n_15455;
and3_13902: n_15451 <=  n_15452  AND n_15453  AND n_15454;
delay_13903: n_15452  <= TRANSPORT a_SCH3MODEREG_F4_G  ;
delay_13904: n_15453  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
delay_13905: n_15454  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and3_13906: n_15455 <=  n_15456  AND n_15457  AND n_15458;
delay_13907: n_15456  <= TRANSPORT a_SCH0MODEREG_F4_G  ;
inv_13908: n_15457  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
inv_13909: n_15458  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and1_13910: n_15459 <=  gnd;
delay_13911: a_N1742_aNOT  <= TRANSPORT a_EQ501  ;
xor2_13912: a_EQ501 <=  n_15462  XOR n_15469;
or2_13913: n_15462 <=  n_15463  OR n_15466;
and2_13914: n_15463 <=  n_15464  AND n_15465;
delay_13915: n_15464  <= TRANSPORT a_N66  ;
delay_13916: n_15465  <= TRANSPORT a_LC8_E2  ;
and2_13917: n_15466 <=  n_15467  AND n_15468;
delay_13918: n_15467  <= TRANSPORT a_N66  ;
delay_13919: n_15468  <= TRANSPORT a_LC7_E2  ;
and1_13920: n_15469 <=  gnd;
delay_13921: a_LC4_E23  <= TRANSPORT a_EQ057  ;
xor2_13922: a_EQ057 <=  n_15472  XOR n_15480;
or3_13923: n_15472 <=  n_15473  OR n_15475  OR n_15477;
and1_13924: n_15473 <=  n_15474;
delay_13925: n_15474  <= TRANSPORT a_LC3_E18  ;
and1_13926: n_15475 <=  n_15476;
delay_13927: n_15476  <= TRANSPORT a_N1742_aNOT  ;
and2_13928: n_15477 <=  n_15478  AND n_15479;
delay_13929: n_15478  <= TRANSPORT a_STEMPORARYREG_F6_G  ;
delay_13930: n_15479  <= TRANSPORT a_N1830  ;
and1_13931: n_15480 <=  gnd;
delay_13932: a_LC3_E23  <= TRANSPORT a_EQ058  ;
xor2_13933: a_EQ058 <=  n_15483  XOR n_15493;
or3_13934: n_15483 <=  n_15484  OR n_15487  OR n_15490;
and2_13935: n_15484 <=  n_15485  AND n_15486;
delay_13936: n_15485  <= TRANSPORT a_N1584  ;
delay_13937: n_15486  <= TRANSPORT a_STEMPORARYREG_F6_G  ;
and2_13938: n_15487 <=  n_15488  AND n_15489;
inv_13939: n_15488  <= TRANSPORT NOT a_N1584  ;
delay_13940: n_15489  <= TRANSPORT a_SADDRESSOUT_F14_G  ;
and2_13941: n_15490 <=  n_15491  AND n_15492;
inv_13942: n_15491  <= TRANSPORT NOT a_N2563_aNOT  ;
delay_13943: n_15492  <= TRANSPORT a_SADDRESSOUT_F14_G  ;
and1_13944: n_15493 <=  gnd;
delay_13945: a_G142  <= TRANSPORT a_EQ059  ;
xor2_13946: a_EQ059 <=  n_15495  XOR n_15508;
or4_13947: n_15495 <=  n_15496  OR n_15499  OR n_15502  OR n_15505;
and2_13948: n_15496 <=  n_15497  AND n_15498;
delay_13949: n_15497  <= TRANSPORT a_LC4_E23  ;
delay_13950: n_15498  <= TRANSPORT a_LC3_E23  ;
and2_13951: n_15499 <=  n_15500  AND n_15501;
delay_13952: n_15500  <= TRANSPORT a_SAEN_aNOT  ;
delay_13953: n_15501  <= TRANSPORT a_LC4_E23  ;
and2_13954: n_15502 <=  n_15503  AND n_15504;
delay_13955: n_15503  <= TRANSPORT a_LC5_B7  ;
delay_13956: n_15504  <= TRANSPORT a_LC3_E23  ;
and2_13957: n_15505 <=  n_15506  AND n_15507;
delay_13958: n_15506  <= TRANSPORT a_SAEN_aNOT  ;
delay_13959: n_15507  <= TRANSPORT a_LC5_B7  ;
and1_13960: n_15508 <=  gnd;
delay_13961: a_N565_aNOT  <= TRANSPORT a_EQ269  ;
xor2_13962: a_EQ269 <=  n_15511  XOR n_15520;
or2_13963: n_15511 <=  n_15512  OR n_15516;
and3_13964: n_15512 <=  n_15513  AND n_15514  AND n_15515;
inv_13965: n_15513  <= TRANSPORT NOT a_N2367  ;
inv_13966: n_15514  <= TRANSPORT NOT a_SCOMMANDREG_F6_G  ;
delay_13967: n_15515  <= TRANSPORT a_N4182  ;
and3_13968: n_15516 <=  n_15517  AND n_15518  AND n_15519;
inv_13969: n_15517  <= TRANSPORT NOT a_N2367  ;
delay_13970: n_15518  <= TRANSPORT a_SCOMMANDREG_F6_G  ;
inv_13971: n_15519  <= TRANSPORT NOT a_N4182  ;
and1_13972: n_15520 <=  gnd;
delay_13973: a_LC8_D15  <= TRANSPORT a_EQ161  ;
xor2_13974: a_EQ161 <=  n_15523  XOR n_15530;
or2_13975: n_15523 <=  n_15524  OR n_15527;
and2_13976: n_15524 <=  n_15525  AND n_15526;
inv_13977: n_15525  <= TRANSPORT NOT a_N77_aNOT  ;
delay_13978: n_15526  <= TRANSPORT a_SCH2ADDRREG_F7_G  ;
and2_13979: n_15527 <=  n_15528  AND n_15529;
inv_13980: n_15528  <= TRANSPORT NOT a_N2347  ;
delay_13981: n_15529  <= TRANSPORT a_SCH3WRDCNTREG_F7_G  ;
and1_13982: n_15530 <=  gnd;
delay_13983: a_LC7_D15  <= TRANSPORT a_EQ162  ;
xor2_13984: a_EQ162 <=  n_15533  XOR n_15540;
or2_13985: n_15533 <=  n_15534  OR n_15537;
and2_13986: n_15534 <=  n_15535  AND n_15536;
inv_13987: n_15535  <= TRANSPORT NOT a_N62_aNOT  ;
delay_13988: n_15536  <= TRANSPORT a_SCH2WRDCNTREG_F7_G  ;
and2_13989: n_15537 <=  n_15538  AND n_15539;
inv_13990: n_15538  <= TRANSPORT NOT a_N2351  ;
delay_13991: n_15539  <= TRANSPORT a_SCH1WRDCNTREG_F7_G  ;
and1_13992: n_15540 <=  gnd;
delay_13993: a_LC6_D15  <= TRANSPORT a_EQ163  ;
xor2_13994: a_EQ163 <=  n_15543  XOR n_15550;
or2_13995: n_15543 <=  n_15544  OR n_15547;
and2_13996: n_15544 <=  n_15545  AND n_15546;
delay_13997: n_15545  <= TRANSPORT a_N2354_aNOT  ;
delay_13998: n_15546  <= TRANSPORT a_SCH0ADDRREG_F7_G  ;
and2_13999: n_15547 <=  n_15548  AND n_15549;
inv_14000: n_15548  <= TRANSPORT NOT a_N2348  ;
delay_14001: n_15549  <= TRANSPORT a_SCH3ADDRREG_F7_G  ;
and1_14002: n_15550 <=  gnd;
delay_14003: a_LC5_D15  <= TRANSPORT a_EQ164  ;
xor2_14004: a_EQ164 <=  n_15553  XOR n_15560;
or2_14005: n_15553 <=  n_15554  OR n_15557;
and2_14006: n_15554 <=  n_15555  AND n_15556;
inv_14007: n_15555  <= TRANSPORT NOT a_N2352  ;
delay_14008: n_15556  <= TRANSPORT a_SCH1ADDRREG_F7_G  ;
and2_14009: n_15557 <=  n_15558  AND n_15559;
inv_14010: n_15558  <= TRANSPORT NOT a_N2353  ;
delay_14011: n_15559  <= TRANSPORT a_SCH0WRDCNTREG_F7_G  ;
and1_14012: n_15560 <=  gnd;
delay_14013: a_LC3_D15  <= TRANSPORT a_EQ165  ;
xor2_14014: a_EQ165 <=  n_15563  XOR n_15572;
or4_14015: n_15563 <=  n_15564  OR n_15566  OR n_15568  OR n_15570;
and1_14016: n_15564 <=  n_15565;
delay_14017: n_15565  <= TRANSPORT a_LC8_D15  ;
and1_14018: n_15566 <=  n_15567;
delay_14019: n_15567  <= TRANSPORT a_LC7_D15  ;
and1_14020: n_15568 <=  n_15569;
delay_14021: n_15569  <= TRANSPORT a_LC6_D15  ;
and1_14022: n_15570 <=  n_15571;
delay_14023: n_15571  <= TRANSPORT a_LC5_D15  ;
and1_14024: n_15572 <=  gnd;
delay_14025: a_LC6_D13  <= TRANSPORT a_EQ166  ;
xor2_14026: a_EQ166 <=  n_15575  XOR n_15582;
or2_14027: n_15575 <=  n_15576  OR n_15579;
and2_14028: n_15576 <=  n_15577  AND n_15578;
inv_14029: n_15577  <= TRANSPORT NOT a_N77_aNOT  ;
delay_14030: n_15578  <= TRANSPORT a_SCH2ADDRREG_F15_G  ;
and2_14031: n_15579 <=  n_15580  AND n_15581;
inv_14032: n_15580  <= TRANSPORT NOT a_N2347  ;
delay_14033: n_15581  <= TRANSPORT a_SH3WRDCNTREG_F15_G  ;
and1_14034: n_15582 <=  gnd;
delay_14035: a_LC5_D13  <= TRANSPORT a_EQ167  ;
xor2_14036: a_EQ167 <=  n_15585  XOR n_15592;
or2_14037: n_15585 <=  n_15586  OR n_15589;
and2_14038: n_15586 <=  n_15587  AND n_15588;
inv_14039: n_15587  <= TRANSPORT NOT a_N62_aNOT  ;
delay_14040: n_15588  <= TRANSPORT a_SH2WRDCNTREG_F15_G  ;
and2_14041: n_15589 <=  n_15590  AND n_15591;
inv_14042: n_15590  <= TRANSPORT NOT a_N2351  ;
delay_14043: n_15591  <= TRANSPORT a_SH1WRDCNTREG_F15_G  ;
and1_14044: n_15592 <=  gnd;
delay_14045: a_LC4_D13  <= TRANSPORT a_EQ168  ;
xor2_14046: a_EQ168 <=  n_15595  XOR n_15602;
or2_14047: n_15595 <=  n_15596  OR n_15599;
and2_14048: n_15596 <=  n_15597  AND n_15598;
delay_14049: n_15597  <= TRANSPORT a_N2354_aNOT  ;
delay_14050: n_15598  <= TRANSPORT a_SCH0ADDRREG_F15_G  ;
and2_14051: n_15599 <=  n_15600  AND n_15601;
inv_14052: n_15600  <= TRANSPORT NOT a_N2348  ;
delay_14053: n_15601  <= TRANSPORT a_SCH3ADDRREG_F15_G  ;
and1_14054: n_15602 <=  gnd;
delay_14055: a_LC2_D13  <= TRANSPORT a_EQ169  ;
xor2_14056: a_EQ169 <=  n_15605  XOR n_15612;
or2_14057: n_15605 <=  n_15606  OR n_15609;
and2_14058: n_15606 <=  n_15607  AND n_15608;
inv_14059: n_15607  <= TRANSPORT NOT a_N2352  ;
delay_14060: n_15608  <= TRANSPORT a_SCH1ADDRREG_F15_G  ;
and2_14061: n_15609 <=  n_15610  AND n_15611;
inv_14062: n_15610  <= TRANSPORT NOT a_N2353  ;
delay_14063: n_15611  <= TRANSPORT a_SH0WRDCNTREG_F15_G  ;
and1_14064: n_15612 <=  gnd;
delay_14065: a_LC1_D13  <= TRANSPORT a_EQ170  ;
xor2_14066: a_EQ170 <=  n_15615  XOR n_15624;
or4_14067: n_15615 <=  n_15616  OR n_15618  OR n_15620  OR n_15622;
and1_14068: n_15616 <=  n_15617;
delay_14069: n_15617  <= TRANSPORT a_LC6_D13  ;
and1_14070: n_15618 <=  n_15619;
delay_14071: n_15619  <= TRANSPORT a_LC5_D13  ;
and1_14072: n_15620 <=  n_15621;
delay_14073: n_15621  <= TRANSPORT a_LC4_D13  ;
and1_14074: n_15622 <=  n_15623;
delay_14075: n_15623  <= TRANSPORT a_LC2_D13  ;
and1_14076: n_15624 <=  gnd;
delay_14077: a_LC3_D13  <= TRANSPORT a_EQ171  ;
xor2_14078: a_EQ171 <=  n_15627  XOR n_15636;
or3_14079: n_15627 <=  n_15628  OR n_15630  OR n_15633;
and1_14080: n_15628 <=  n_15629;
delay_14081: n_15629  <= TRANSPORT a_N565_aNOT  ;
and2_14082: n_15630 <=  n_15631  AND n_15632;
inv_14083: n_15631  <= TRANSPORT NOT bytepointer  ;
delay_14084: n_15632  <= TRANSPORT a_LC3_D15  ;
and2_14085: n_15633 <=  n_15634  AND n_15635;
delay_14086: n_15634  <= TRANSPORT bytepointer  ;
delay_14087: n_15635  <= TRANSPORT a_LC1_D13  ;
and1_14088: n_15636 <=  gnd;
delay_14089: a_N1226_aNOT  <= TRANSPORT a_N1226_aNOT_aIN  ;
xor2_14090: a_N1226_aNOT_aIN <=  n_15639  XOR n_15643;
or1_14091: n_15639 <=  n_15640;
and2_14092: n_15640 <=  n_15641  AND n_15642;
inv_14093: n_15641  <= TRANSPORT NOT a_N2557  ;
delay_14094: n_15642  <= TRANSPORT a_SADDRESSOUT_F15_G  ;
and1_14095: n_15643 <=  gnd;
delay_14096: a_LC6_E24  <= TRANSPORT a_EQ160  ;
xor2_14097: a_EQ160 <=  n_15646  XOR n_15654;
or3_14098: n_15646 <=  n_15647  OR n_15649  OR n_15652;
and1_14099: n_15647 <=  n_15648;
delay_14100: n_15648  <= TRANSPORT a_N1226_aNOT  ;
and2_14101: n_15649 <=  n_15650  AND n_15651;
delay_14102: n_15650  <= TRANSPORT a_N1584  ;
delay_14103: n_15651  <= TRANSPORT a_STEMPORARYREG_F7_G  ;
and1_14104: n_15652 <=  n_15653;
delay_14105: n_15653  <= TRANSPORT a_SAEN_aNOT  ;
and1_14106: n_15654 <=  gnd;
delay_14107: a_LC2_E24  <= TRANSPORT a_EQ172  ;
xor2_14108: a_EQ172 <=  n_15657  XOR n_15664;
or2_14109: n_15657 <=  n_15658  OR n_15661;
and2_14110: n_15658 <=  n_15659  AND n_15660;
delay_14111: n_15659  <= TRANSPORT a_STEMPORARYREG_F7_G  ;
delay_14112: n_15660  <= TRANSPORT a_N1830  ;
and2_14113: n_15661 <=  n_15662  AND n_15663;
delay_14114: n_15662  <= TRANSPORT a_N73  ;
delay_14115: n_15663  <= TRANSPORT a_SCOMMANDREG_F7_G  ;
and1_14116: n_15664 <=  gnd;
delay_14117: a_LC7_E15  <= TRANSPORT a_EQ387  ;
xor2_14118: a_EQ387 <=  n_15667  XOR n_15676;
or2_14119: n_15667 <=  n_15668  OR n_15672;
and3_14120: n_15668 <=  n_15669  AND n_15670  AND n_15671;
delay_14121: n_15669  <= TRANSPORT a_SCH3MODEREG_F5_G  ;
delay_14122: n_15670  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
delay_14123: n_15671  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and3_14124: n_15672 <=  n_15673  AND n_15674  AND n_15675;
delay_14125: n_15673  <= TRANSPORT a_SCH1MODEREG_F5_G  ;
inv_14126: n_15674  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
delay_14127: n_15675  <= TRANSPORT a_SMODECOUNTER_F0_G  ;
and1_14128: n_15676 <=  gnd;
delay_14129: a_LC3_E26  <= TRANSPORT a_EQ388  ;
xor2_14130: a_EQ388 <=  n_15679  XOR n_15688;
or2_14131: n_15679 <=  n_15680  OR n_15684;
and3_14132: n_15680 <=  n_15681  AND n_15682  AND n_15683;
delay_14133: n_15681  <= TRANSPORT a_SCH2MODEREG_F5_G  ;
delay_14134: n_15682  <= TRANSPORT a_SMODECOUNTER_F1_G  ;
inv_14135: n_15683  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
and3_14136: n_15684 <=  n_15685  AND n_15686  AND n_15687;
inv_14137: n_15685  <= TRANSPORT NOT a_SMODECOUNTER_F1_G  ;
inv_14138: n_15686  <= TRANSPORT NOT a_SMODECOUNTER_F0_G  ;
delay_14139: n_15687  <= TRANSPORT a_SCH0MODEREG_F5_G  ;
and1_14140: n_15688 <=  gnd;
delay_14141: a_LC1_E24  <= TRANSPORT a_EQ173  ;
xor2_14142: a_EQ173 <=  n_15691  XOR n_15700;
or3_14143: n_15691 <=  n_15692  OR n_15694  OR n_15697;
and1_14144: n_15692 <=  n_15693;
delay_14145: n_15693  <= TRANSPORT a_LC2_E24  ;
and2_14146: n_15694 <=  n_15695  AND n_15696;
delay_14147: n_15695  <= TRANSPORT a_N66  ;
delay_14148: n_15696  <= TRANSPORT a_LC7_E15  ;
and2_14149: n_15697 <=  n_15698  AND n_15699;
delay_14150: n_15698  <= TRANSPORT a_N66  ;
delay_14151: n_15699  <= TRANSPORT a_LC3_E26  ;
and1_14152: n_15700 <=  gnd;
delay_14153: a_G1389  <= TRANSPORT a_EQ174  ;
xor2_14154: a_EQ174 <=  n_15702  XOR n_15712;
or3_14155: n_15702 <=  n_15703  OR n_15706  OR n_15709;
and2_14156: n_15703 <=  n_15704  AND n_15705;
delay_14157: n_15704  <= TRANSPORT a_LC3_D13  ;
delay_14158: n_15705  <= TRANSPORT a_LC6_E24  ;
and2_14159: n_15706 <=  n_15707  AND n_15708;
delay_14160: n_15707  <= TRANSPORT a_LC6_E24  ;
delay_14161: n_15708  <= TRANSPORT a_LC1_E24  ;
and2_14162: n_15709 <=  n_15710  AND n_15711;
delay_14163: n_15710  <= TRANSPORT a_LC5_B7  ;
delay_14164: n_15711  <= TRANSPORT a_LC6_E24  ;
and1_14165: n_15712 <=  gnd;
delay_14166: a_N2588  <= TRANSPORT a_EQ641  ;
xor2_14167: a_EQ641 <=  n_15715  XOR n_15725;
or3_14168: n_15715 <=  n_15716  OR n_15719  OR n_15722;
and2_14169: n_15716 <=  n_15717  AND n_15718;
delay_14170: n_15717  <= TRANSPORT a_N2563_aNOT  ;
inv_14171: n_15718  <= TRANSPORT NOT a_N2358  ;
and2_14172: n_15719 <=  n_15720  AND n_15721;
delay_14173: n_15720  <= TRANSPORT a_N2563_aNOT  ;
inv_14174: n_15721  <= TRANSPORT NOT a_N68_aNOT  ;
and2_14175: n_15722 <=  n_15723  AND n_15724;
delay_14176: n_15723  <= TRANSPORT a_N2563_aNOT  ;
inv_14177: n_15724  <= TRANSPORT NOT a_N1592  ;
and1_14178: n_15725 <=  gnd;
delay_14179: a_G503  <= TRANSPORT a_EQ094  ;
xor2_14180: a_EQ094 <=  n_15727  XOR n_15742;
or4_14181: n_15727 <=  n_15728  OR n_15731  OR n_15734  OR n_15737;
and2_14182: n_15728 <=  n_15729  AND n_15730;
inv_14183: n_15729  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14184: n_15730  <= TRANSPORT NOT a_N2588  ;
and2_14185: n_15731 <=  n_15732  AND n_15733;
inv_14186: n_15732  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
delay_14187: n_15733  <= TRANSPORT a_SCHANNEL_F1_G  ;
and2_14188: n_15734 <=  n_15735  AND n_15736;
inv_14189: n_15735  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
delay_14190: n_15736  <= TRANSPORT a_SCHANNEL_F0_G  ;
and4_14191: n_15737 <=  n_15738  AND n_15739  AND n_15740  AND n_15741;
delay_14192: n_15738  <= TRANSPORT a_SCOMMANDREG_F7_G  ;
inv_14193: n_15739  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
inv_14194: n_15740  <= TRANSPORT NOT a_SCHANNEL_F0_G  ;
delay_14195: n_15741  <= TRANSPORT a_N2588  ;
and1_14196: n_15742 <=  gnd;
delay_14197: a_G502  <= TRANSPORT a_EQ093  ;
xor2_14198: a_EQ093 <=  n_15744  XOR n_15759;
or4_14199: n_15744 <=  n_15745  OR n_15748  OR n_15751  OR n_15754;
and2_14200: n_15745 <=  n_15746  AND n_15747;
inv_14201: n_15746  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
delay_14202: n_15747  <= TRANSPORT a_SCHANNEL_F1_G  ;
and2_14203: n_15748 <=  n_15749  AND n_15750;
inv_14204: n_15749  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14205: n_15750  <= TRANSPORT NOT a_SCHANNEL_F0_G  ;
and2_14206: n_15751 <=  n_15752  AND n_15753;
inv_14207: n_15752  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14208: n_15753  <= TRANSPORT NOT a_N2588  ;
and4_14209: n_15754 <=  n_15755  AND n_15756  AND n_15757  AND n_15758;
delay_14210: n_15755  <= TRANSPORT a_SCOMMANDREG_F7_G  ;
inv_14211: n_15756  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
delay_14212: n_15757  <= TRANSPORT a_SCHANNEL_F0_G  ;
delay_14213: n_15758  <= TRANSPORT a_N2588  ;
and1_14214: n_15759 <=  gnd;
delay_14215: a_G1464  <= TRANSPORT a_EQ176  ;
xor2_14216: a_EQ176 <=  n_15761  XOR n_15776;
or4_14217: n_15761 <=  n_15762  OR n_15765  OR n_15768  OR n_15771;
and2_14218: n_15762 <=  n_15763  AND n_15764;
inv_14219: n_15763  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14220: n_15764  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and2_14221: n_15765 <=  n_15766  AND n_15767;
inv_14222: n_15766  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
delay_14223: n_15767  <= TRANSPORT a_SCHANNEL_F0_G  ;
and2_14224: n_15768 <=  n_15769  AND n_15770;
inv_14225: n_15769  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14226: n_15770  <= TRANSPORT NOT a_N2588  ;
and4_14227: n_15771 <=  n_15772  AND n_15773  AND n_15774  AND n_15775;
delay_14228: n_15772  <= TRANSPORT a_SCOMMANDREG_F7_G  ;
delay_14229: n_15773  <= TRANSPORT a_SCHANNEL_F1_G  ;
inv_14230: n_15774  <= TRANSPORT NOT a_SCHANNEL_F0_G  ;
delay_14231: n_15775  <= TRANSPORT a_N2588  ;
and1_14232: n_15776 <=  gnd;
delay_14233: a_G1463  <= TRANSPORT a_EQ175  ;
xor2_14234: a_EQ175 <=  n_15778  XOR n_15793;
or4_14235: n_15778 <=  n_15779  OR n_15782  OR n_15785  OR n_15788;
and2_14236: n_15779 <=  n_15780  AND n_15781;
inv_14237: n_15780  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14238: n_15781  <= TRANSPORT NOT a_SCHANNEL_F1_G  ;
and2_14239: n_15782 <=  n_15783  AND n_15784;
inv_14240: n_15783  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14241: n_15784  <= TRANSPORT NOT a_SCHANNEL_F0_G  ;
and2_14242: n_15785 <=  n_15786  AND n_15787;
inv_14243: n_15786  <= TRANSPORT NOT a_SCOMMANDREG_F7_G  ;
inv_14244: n_15787  <= TRANSPORT NOT a_N2588  ;
and4_14245: n_15788 <=  n_15789  AND n_15790  AND n_15791  AND n_15792;
delay_14246: n_15789  <= TRANSPORT a_SCOMMANDREG_F7_G  ;
delay_14247: n_15790  <= TRANSPORT a_SCHANNEL_F1_G  ;
delay_14248: n_15791  <= TRANSPORT a_SCHANNEL_F0_G  ;
delay_14249: n_15792  <= TRANSPORT a_N2588  ;
and1_14250: n_15793 <=  gnd;
delay_14251: a_N2400  <= TRANSPORT a_EQ578  ;
xor2_14252: a_EQ578 <=  n_15796  XOR n_15805;
or4_14253: n_15796 <=  n_15797  OR n_15799  OR n_15801  OR n_15803;
and1_14254: n_15797 <=  n_15798;
inv_14255: n_15798  <= TRANSPORT NOT a_N2358  ;
and1_14256: n_15799 <=  n_15800;
inv_14257: n_15800  <= TRANSPORT NOT a_N1566  ;
and1_14258: n_15801 <=  n_15802;
inv_14259: n_15802  <= TRANSPORT NOT a_LC4_B25_aNOT  ;
and1_14260: n_15803 <=  n_15804;
delay_14261: n_15804  <= TRANSPORT a_N2372_aNOT  ;
and1_14262: n_15805 <=  gnd;
delay_14263: a_LC5_B5  <= TRANSPORT a_EQ1172  ;
xor2_14264: a_EQ1172 <=  n_15808  XOR n_15815;
or3_14265: n_15808 <=  n_15809  OR n_15811  OR n_15813;
and1_14266: n_15809 <=  n_15810;
delay_14267: n_15810  <= TRANSPORT a_N2400  ;
and1_14268: n_15811 <=  n_15812;
delay_14269: n_15812  <= TRANSPORT a_N70  ;
and1_14270: n_15813 <=  n_15814;
inv_14271: n_15814  <= TRANSPORT NOT a_N2563_aNOT  ;
and1_14272: n_15815 <=  gnd;
delay_14273: a_N2368  <= TRANSPORT a_EQ564  ;
xor2_14274: a_EQ564 <=  n_15818  XOR n_15826;
or3_14275: n_15818 <=  n_15819  OR n_15822  OR n_15824;
and2_14276: n_15819 <=  n_15820  AND n_15821;
delay_14277: n_15820  <= TRANSPORT a_LC6_E22  ;
delay_14278: n_15821  <= TRANSPORT a_LC5_E22  ;
and1_14279: n_15822 <=  n_15823;
delay_14280: n_15823  <= TRANSPORT a_LC4_E22  ;
and1_14281: n_15824 <=  n_15825;
delay_14282: n_15825  <= TRANSPORT a_LC6_E10  ;
and1_14283: n_15826 <=  gnd;
delay_14284: a_LC7_B5  <= TRANSPORT a_EQ1171  ;
xor2_14285: a_EQ1171 <=  n_15829  XOR n_15837;
or2_14286: n_15829 <=  n_15830  OR n_15834;
and3_14287: n_15830 <=  n_15831  AND n_15832  AND n_15833;
inv_14288: n_15831  <= TRANSPORT NOT a_LC1_B23_aNOT  ;
inv_14289: n_15832  <= TRANSPORT NOT a_N820  ;
delay_14290: n_15833  <= TRANSPORT a_N2368  ;
and2_14291: n_15834 <=  n_15835  AND n_15836;
inv_14292: n_15835  <= TRANSPORT NOT a_N67_aNOT  ;
delay_14293: n_15836  <= TRANSPORT a_N2368  ;
and1_14294: n_15837 <=  gnd;
delay_14295: a_LC2_B5  <= TRANSPORT a_EQ447  ;
xor2_14296: a_EQ447 <=  n_15840  XOR n_15850;
or3_14297: n_15840 <=  n_15841  OR n_15844  OR n_15847;
and2_14298: n_15841 <=  n_15842  AND n_15843;
delay_14299: n_15842  <= TRANSPORT a_N1467  ;
inv_14300: n_15843  <= TRANSPORT NOT a_N823  ;
and2_14301: n_15844 <=  n_15845  AND n_15846;
delay_14302: n_15845  <= TRANSPORT a_N1467  ;
delay_14303: n_15846  <= TRANSPORT a_N822  ;
and2_14304: n_15847 <=  n_15848  AND n_15849;
delay_14305: n_15848  <= TRANSPORT a_N1467  ;
inv_14306: n_15849  <= TRANSPORT NOT a_SCOMMANDREG_F5_G  ;
and1_14307: n_15850 <=  gnd;
delay_14308: a_N1468  <= TRANSPORT a_EQ449  ;
xor2_14309: a_EQ449 <=  n_15853  XOR n_15862;
or3_14310: n_15853 <=  n_15854  OR n_15857  OR n_15860;
and2_14311: n_15854 <=  n_15855  AND n_15856;
inv_14312: n_15855  <= TRANSPORT NOT a_N823  ;
delay_14313: n_15856  <= TRANSPORT a_N2368  ;
and2_14314: n_15857 <=  n_15858  AND n_15859;
inv_14315: n_15858  <= TRANSPORT NOT a_SCOMMANDREG_F5_G  ;
inv_14316: n_15859  <= TRANSPORT NOT a_N823  ;
and1_14317: n_15860 <=  n_15861;
delay_14318: n_15861  <= TRANSPORT a_N820  ;
and1_14319: n_15862 <=  gnd;
delay_14320: a_SNMEMW  <= TRANSPORT a_EQ1170  ;
xor2_14321: a_EQ1170 <=  n_15864  XOR n_15872;
or3_14322: n_15864 <=  n_15865  OR n_15867  OR n_15869;
and1_14323: n_15865 <=  n_15866;
delay_14324: n_15866  <= TRANSPORT a_LC5_B5  ;
and1_14325: n_15867 <=  n_15868;
delay_14326: n_15868  <= TRANSPORT a_LC7_B5  ;
and2_14327: n_15869 <=  n_15870  AND n_15871;
delay_14328: n_15870  <= TRANSPORT a_LC2_B5  ;
delay_14329: n_15871  <= TRANSPORT a_N1468  ;
and1_14330: n_15872 <=  gnd;
delay_14331: a_LC5_B25  <= TRANSPORT a_EQ1168  ;
xor2_14332: a_EQ1168 <=  n_15875  XOR n_15884;
or4_14333: n_15875 <=  n_15876  OR n_15878  OR n_15880  OR n_15882;
and1_14334: n_15876 <=  n_15877;
inv_14335: n_15877  <= TRANSPORT NOT a_LC4_B25_aNOT  ;
and1_14336: n_15878 <=  n_15879;
inv_14337: n_15879  <= TRANSPORT NOT a_N2374  ;
and1_14338: n_15880 <=  n_15881;
delay_14339: n_15881  <= TRANSPORT a_N2372_aNOT  ;
and1_14340: n_15882 <=  n_15883;
delay_14341: n_15883  <= TRANSPORT a_N70  ;
and1_14342: n_15884 <=  gnd;
delay_14343: a_SNIOWOUT  <= TRANSPORT a_EQ1167  ;
xor2_14344: a_EQ1167 <=  n_15886  XOR n_15894;
or3_14345: n_15886 <=  n_15887  OR n_15889  OR n_15892;
and1_14346: n_15887 <=  n_15888;
delay_14347: n_15888  <= TRANSPORT a_LC5_B25  ;
and2_14348: n_15889 <=  n_15890  AND n_15891;
inv_14349: n_15890  <= TRANSPORT NOT a_N2356  ;
inv_14350: n_15891  <= TRANSPORT NOT a_SCOMMANDREG_F5_G  ;
and1_14351: n_15892 <=  n_15893;
inv_14352: n_15893  <= TRANSPORT NOT a_N1580_aNOT  ;
and1_14353: n_15894 <=  gnd;
delay_14354: a_LC2_B20  <= TRANSPORT a_EQ1166  ;
xor2_14355: a_EQ1166 <=  n_15897  XOR n_15906;
or4_14356: n_15897 <=  n_15898  OR n_15900  OR n_15902  OR n_15904;
and1_14357: n_15898 <=  n_15899;
delay_14358: n_15899  <= TRANSPORT a_N70  ;
and1_14359: n_15900 <=  n_15901;
inv_14360: n_15901  <= TRANSPORT NOT a_N71_aNOT  ;
and1_14361: n_15902 <=  n_15903;
inv_14362: n_15903  <= TRANSPORT NOT a_N2374  ;
and1_14363: n_15904 <=  n_15905;
delay_14364: n_15905  <= TRANSPORT a_N2400  ;
and1_14365: n_15906 <=  gnd;
delay_14366: a_SNIOROUT  <= TRANSPORT a_EQ1165  ;
xor2_14367: a_EQ1165 <=  n_15908  XOR n_15916;
or3_14368: n_15908 <=  n_15909  OR n_15911  OR n_15914;
and1_14369: n_15909 <=  n_15910;
delay_14370: n_15910  <= TRANSPORT a_LC2_B20  ;
and2_14371: n_15911 <=  n_15912  AND n_15913;
inv_14372: n_15912  <= TRANSPORT NOT a_N1592  ;
delay_14373: n_15913  <= TRANSPORT a_N2368  ;
and1_14374: n_15914 <=  n_15915;
inv_14375: n_15915  <= TRANSPORT NOT a_LC8_B20  ;
and1_14376: n_15916 <=  gnd;
delay_14377: a_N1252  <= TRANSPORT a_EQ396  ;
xor2_14378: a_EQ396 <=  n_15919  XOR n_15934;
or4_14379: n_15919 <=  n_15920  OR n_15924  OR n_15927  OR n_15931;
and3_14380: n_15920 <=  n_15921  AND n_15922  AND n_15923;
delay_14381: n_15921  <= TRANSPORT a_N820  ;
inv_14382: n_15922  <= TRANSPORT NOT a_N822  ;
inv_14383: n_15923  <= TRANSPORT NOT a_N823  ;
and2_14384: n_15924 <=  n_15925  AND n_15926;
delay_14385: n_15925  <= TRANSPORT a_N820  ;
delay_14386: n_15926  <= TRANSPORT a_N821  ;
and3_14387: n_15927 <=  n_15928  AND n_15929  AND n_15930;
inv_14388: n_15928  <= TRANSPORT NOT a_N820  ;
delay_14389: n_15929  <= TRANSPORT a_N822  ;
inv_14390: n_15930  <= TRANSPORT NOT a_N821  ;
and2_14391: n_15931 <=  n_15932  AND n_15933;
delay_14392: n_15932  <= TRANSPORT a_N822  ;
delay_14393: n_15933  <= TRANSPORT a_N823  ;
and1_14394: n_15934 <=  gnd;
delay_14395: a_SDBEN  <= TRANSPORT a_EQ1131  ;
xor2_14396: a_EQ1131 <=  n_15936  XOR n_15943;
or2_14397: n_15936 <=  n_15937  OR n_15940;
and2_14398: n_15937 <=  n_15938  AND n_15939;
inv_14399: n_15938  <= TRANSPORT NOT niorin  ;
inv_14400: n_15939  <= TRANSPORT NOT ncs  ;
and2_14401: n_15940 <=  n_15941  AND n_15942;
delay_14402: n_15941  <= TRANSPORT a_N2563_aNOT  ;
delay_14403: n_15942  <= TRANSPORT a_N1252  ;
and1_14404: n_15943 <=  gnd;
delay_14405: a_LC6_B16_aNOT  <= TRANSPORT a_LC6_B16_aNOT_aIN  ;
xor2_14406: a_LC6_B16_aNOT_aIN <=  n_15945  XOR n_15950;
or2_14407: n_15945 <=  n_15946  OR n_15948;
and1_14408: n_15946 <=  n_15947;
inv_14409: n_15947  <= TRANSPORT NOT a_N2563_aNOT  ;
and1_14410: n_15948 <=  n_15949;
inv_14411: n_15949  <= TRANSPORT NOT a_N1566  ;
and1_14412: n_15950 <=  gnd;
delay_14413: a_N2370_aNOT  <= TRANSPORT a_N2370_aNOT_aIN  ;
xor2_14414: a_N2370_aNOT_aIN <=  n_15953  XOR n_15958;
or1_14415: n_15953 <=  n_15954;
and3_14416: n_15954 <=  n_15955  AND n_15956  AND n_15957;
delay_14417: n_15955  <= TRANSPORT a_N822  ;
delay_14418: n_15956  <= TRANSPORT a_N821  ;
delay_14419: n_15957  <= TRANSPORT a_N823  ;
and1_14420: n_15958 <=  gnd;
delay_14421: a_SADSTB  <= TRANSPORT a_EQ862  ;
xor2_14422: a_EQ862 <=  n_15960  XOR n_15970;
or3_14423: n_15960 <=  n_15961  OR n_15964  OR n_15967;
and2_14424: n_15961 <=  n_15962  AND n_15963;
delay_14425: n_15962  <= TRANSPORT a_N2563_aNOT  ;
delay_14426: n_15963  <= TRANSPORT a_N2370_aNOT  ;
and2_14427: n_15964 <=  n_15965  AND n_15966;
delay_14428: n_15965  <= TRANSPORT a_N2563_aNOT  ;
inv_14429: n_15966  <= TRANSPORT NOT a_N2358  ;
and2_14430: n_15967 <=  n_15968  AND n_15969;
delay_14431: n_15968  <= TRANSPORT a_N2563_aNOT  ;
inv_14432: n_15969  <= TRANSPORT NOT a_N2374  ;
and1_14433: n_15970 <=  gnd;
delay_14434: a_N87  <= TRANSPORT a_EQ196  ;
xor2_14435: a_EQ196 <=  n_15972  XOR n_15977;
or2_14436: n_15972 <=  n_15973  OR n_15975;
and1_14437: n_15973 <=  n_15974;
delay_14438: n_15974  <= TRANSPORT ncs  ;
and1_14439: n_15975 <=  n_15976;
delay_14440: n_15976  <= TRANSPORT niowin  ;
and1_14441: n_15977 <=  gnd;
delay_14442: a_LC6_D6  <= TRANSPORT a_EQ633  ;
xor2_14443: a_EQ633 <=  n_15979  XOR n_15984;
or2_14444: n_15979 <=  n_15980  OR n_15982;
and1_14445: n_15980 <=  n_15981;
delay_14446: n_15981  <= TRANSPORT bytepointer  ;
and1_14447: n_15982 <=  n_15983;
delay_14448: n_15983  <= TRANSPORT a_N87  ;
and1_14449: n_15984 <=  gnd;
delay_14450: a_N2351  <= TRANSPORT a_EQ555  ;
xor2_14451: a_EQ555 <=  n_15986  XOR n_15995;
or4_14452: n_15986 <=  n_15987  OR n_15989  OR n_15991  OR n_15993;
and1_14453: n_15987 <=  n_15988;
inv_14454: n_15988  <= TRANSPORT NOT ain(0)  ;
and1_14455: n_15989 <=  n_15990;
delay_14456: n_15990  <= TRANSPORT ain(3)  ;
and1_14457: n_15991 <=  n_15992;
delay_14458: n_15992  <= TRANSPORT ain(2)  ;
and1_14459: n_15993 <=  n_15994;
inv_14460: n_15994  <= TRANSPORT NOT ain(1)  ;
and1_14461: n_15995 <=  gnd;
delay_14462: a_N2576_aNOT  <= TRANSPORT a_EQ628  ;
xor2_14463: a_EQ628 <=  n_15997  XOR n_16002;
or2_14464: n_15997 <=  n_15998  OR n_16000;
and1_14465: n_15998 <=  n_15999;
delay_14466: n_15999  <= TRANSPORT a_LC6_D6  ;
and1_14467: n_16000 <=  n_16001;
delay_14468: n_16001  <= TRANSPORT a_N2351  ;
and1_14469: n_16002 <=  gnd;
dff_14470: DFF_a8237

    PORT MAP ( D => a_EQ964, CLK => a_SCH1BWORDOUT_F1_G_aCLK, CLRN => a_SCH1BWORDOUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F1_G);
inv_14471: a_SCH1BWORDOUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14472: a_EQ964 <=  n_16009  XOR n_16016;
or2_14473: n_16009 <=  n_16010  OR n_16013;
and2_14474: n_16010 <=  n_16011  AND n_16012;
inv_14475: n_16011  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_14476: n_16012  <= TRANSPORT dbin(1)  ;
and2_14477: n_16013 <=  n_16014  AND n_16015;
delay_14478: n_16014  <= TRANSPORT a_N2576_aNOT  ;
delay_14479: n_16015  <= TRANSPORT a_SCH1BWORDOUT_F1_G  ;
and1_14480: n_16016 <=  gnd;
delay_14481: n_16017  <= TRANSPORT clk  ;
filter_14482: FILTER_a8237

    PORT MAP (IN1 => n_16017, Y => a_SCH1BWORDOUT_F1_G_aCLK);
delay_14483: a_LC3_D22  <= TRANSPORT a_EQ635  ;
xor2_14484: a_EQ635 <=  n_16020  XOR n_16025;
or2_14485: n_16020 <=  n_16021  OR n_16023;
and1_14486: n_16021 <=  n_16022;
inv_14487: n_16022  <= TRANSPORT NOT bytepointer  ;
and1_14488: n_16023 <=  n_16024;
delay_14489: n_16024  <= TRANSPORT a_N87  ;
and1_14490: n_16025 <=  gnd;
delay_14491: a_N2577_aNOT  <= TRANSPORT a_EQ629  ;
xor2_14492: a_EQ629 <=  n_16027  XOR n_16032;
or2_14493: n_16027 <=  n_16028  OR n_16030;
and1_14494: n_16028 <=  n_16029;
delay_14495: n_16029  <= TRANSPORT a_LC3_D22  ;
and1_14496: n_16030 <=  n_16031;
delay_14497: n_16031  <= TRANSPORT a_N2351  ;
and1_14498: n_16032 <=  gnd;
dff_14499: DFF_a8237

    PORT MAP ( D => a_EQ972, CLK => a_SCH1BWORDOUT_F9_G_aCLK, CLRN => a_SCH1BWORDOUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F9_G);
inv_14500: a_SCH1BWORDOUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14501: a_EQ972 <=  n_16039  XOR n_16046;
or2_14502: n_16039 <=  n_16040  OR n_16043;
and2_14503: n_16040 <=  n_16041  AND n_16042;
inv_14504: n_16041  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_14505: n_16042  <= TRANSPORT dbin(1)  ;
and2_14506: n_16043 <=  n_16044  AND n_16045;
delay_14507: n_16044  <= TRANSPORT a_N2577_aNOT  ;
delay_14508: n_16045  <= TRANSPORT a_SCH1BWORDOUT_F9_G  ;
and1_14509: n_16046 <=  gnd;
delay_14510: n_16047  <= TRANSPORT clk  ;
filter_14511: FILTER_a8237

    PORT MAP (IN1 => n_16047, Y => a_SCH1BWORDOUT_F9_G_aCLK);
dff_14512: DFF_a8237

    PORT MAP ( D => a_EQ973, CLK => a_SCH1BWORDOUT_F10_G_aCLK, CLRN => a_SCH1BWORDOUT_F10_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F10_G);
inv_14513: a_SCH1BWORDOUT_F10_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14514: a_EQ973 <=  n_16055  XOR n_16062;
or2_14515: n_16055 <=  n_16056  OR n_16059;
and2_14516: n_16056 <=  n_16057  AND n_16058;
inv_14517: n_16057  <= TRANSPORT NOT a_N2577_aNOT  ;
delay_14518: n_16058  <= TRANSPORT dbin(2)  ;
and2_14519: n_16059 <=  n_16060  AND n_16061;
delay_14520: n_16060  <= TRANSPORT a_N2577_aNOT  ;
delay_14521: n_16061  <= TRANSPORT a_SCH1BWORDOUT_F10_G  ;
and1_14522: n_16062 <=  gnd;
delay_14523: n_16063  <= TRANSPORT clk  ;
filter_14524: FILTER_a8237

    PORT MAP (IN1 => n_16063, Y => a_SCH1BWORDOUT_F10_G_aCLK);
delay_14525: a_N2347  <= TRANSPORT a_EQ553  ;
xor2_14526: a_EQ553 <=  n_16066  XOR n_16075;
or4_14527: n_16066 <=  n_16067  OR n_16069  OR n_16071  OR n_16073;
and1_14528: n_16067 <=  n_16068;
inv_14529: n_16068  <= TRANSPORT NOT ain(0)  ;
and1_14530: n_16069 <=  n_16070;
delay_14531: n_16070  <= TRANSPORT ain(3)  ;
and1_14532: n_16071 <=  n_16072;
inv_14533: n_16072  <= TRANSPORT NOT ain(2)  ;
and1_14534: n_16073 <=  n_16074;
inv_14535: n_16074  <= TRANSPORT NOT ain(1)  ;
and1_14536: n_16075 <=  gnd;
delay_14537: a_N2572_aNOT  <= TRANSPORT a_EQ625  ;
xor2_14538: a_EQ625 <=  n_16077  XOR n_16084;
or3_14539: n_16077 <=  n_16078  OR n_16080  OR n_16082;
and1_14540: n_16078 <=  n_16079;
delay_14541: n_16079  <= TRANSPORT bytepointer  ;
and1_14542: n_16080 <=  n_16081;
delay_14543: n_16081  <= TRANSPORT a_N87  ;
and1_14544: n_16082 <=  n_16083;
delay_14545: n_16083  <= TRANSPORT a_N2347  ;
and1_14546: n_16084 <=  gnd;
dff_14547: DFF_a8237

    PORT MAP ( D => a_EQ1097, CLK => a_SCH3BWORDOUT_F6_G_aCLK, CLRN => a_SCH3BWORDOUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F6_G);
inv_14548: a_SCH3BWORDOUT_F6_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14549: a_EQ1097 <=  n_16091  XOR n_16098;
or2_14550: n_16091 <=  n_16092  OR n_16095;
and2_14551: n_16092 <=  n_16093  AND n_16094;
inv_14552: n_16093  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_14553: n_16094  <= TRANSPORT dbin(6)  ;
and2_14554: n_16095 <=  n_16096  AND n_16097;
delay_14555: n_16096  <= TRANSPORT a_N2572_aNOT  ;
delay_14556: n_16097  <= TRANSPORT a_SCH3BWORDOUT_F6_G  ;
and1_14557: n_16098 <=  gnd;
delay_14558: n_16099  <= TRANSPORT clk  ;
filter_14559: FILTER_a8237

    PORT MAP (IN1 => n_16099, Y => a_SCH3BWORDOUT_F6_G_aCLK);
dff_14560: DFF_a8237

    PORT MAP ( D => a_EQ1092, CLK => a_SCH3BWORDOUT_F1_G_aCLK, CLRN => a_SCH3BWORDOUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH3BWORDOUT_F1_G);
inv_14561: a_SCH3BWORDOUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14562: a_EQ1092 <=  n_16107  XOR n_16114;
or2_14563: n_16107 <=  n_16108  OR n_16111;
and2_14564: n_16108 <=  n_16109  AND n_16110;
inv_14565: n_16109  <= TRANSPORT NOT a_N2572_aNOT  ;
delay_14566: n_16110  <= TRANSPORT dbin(1)  ;
and2_14567: n_16111 <=  n_16112  AND n_16113;
delay_14568: n_16112  <= TRANSPORT a_N2572_aNOT  ;
delay_14569: n_16113  <= TRANSPORT a_SCH3BWORDOUT_F1_G  ;
and1_14570: n_16114 <=  gnd;
delay_14571: n_16115  <= TRANSPORT clk  ;
filter_14572: FILTER_a8237

    PORT MAP (IN1 => n_16115, Y => a_SCH3BWORDOUT_F1_G_aCLK);
delay_14573: a_N62_aNOT  <= TRANSPORT a_EQ183  ;
xor2_14574: a_EQ183 <=  n_16118  XOR n_16127;
or4_14575: n_16118 <=  n_16119  OR n_16121  OR n_16123  OR n_16125;
and1_14576: n_16119 <=  n_16120;
inv_14577: n_16120  <= TRANSPORT NOT ain(0)  ;
and1_14578: n_16121 <=  n_16122;
delay_14579: n_16122  <= TRANSPORT ain(3)  ;
and1_14580: n_16123 <=  n_16124;
inv_14581: n_16124  <= TRANSPORT NOT ain(2)  ;
and1_14582: n_16125 <=  n_16126;
delay_14583: n_16126  <= TRANSPORT ain(1)  ;
and1_14584: n_16127 <=  gnd;
delay_14585: a_N2574_aNOT  <= TRANSPORT a_EQ627  ;
xor2_14586: a_EQ627 <=  n_16129  XOR n_16134;
or2_14587: n_16129 <=  n_16130  OR n_16132;
and1_14588: n_16130 <=  n_16131;
delay_14589: n_16131  <= TRANSPORT a_LC6_D6  ;
and1_14590: n_16132 <=  n_16133;
delay_14591: n_16133  <= TRANSPORT a_N62_aNOT  ;
and1_14592: n_16134 <=  gnd;
dff_14593: DFF_a8237

    PORT MAP ( D => a_EQ1028, CLK => a_SCH2BWORDOUT_F1_G_aCLK, CLRN => a_SCH2BWORDOUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F1_G);
inv_14594: a_SCH2BWORDOUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14595: a_EQ1028 <=  n_16141  XOR n_16148;
or2_14596: n_16141 <=  n_16142  OR n_16145;
and2_14597: n_16142 <=  n_16143  AND n_16144;
inv_14598: n_16143  <= TRANSPORT NOT a_N2574_aNOT  ;
delay_14599: n_16144  <= TRANSPORT dbin(1)  ;
and2_14600: n_16145 <=  n_16146  AND n_16147;
delay_14601: n_16146  <= TRANSPORT a_N2574_aNOT  ;
delay_14602: n_16147  <= TRANSPORT a_SCH2BWORDOUT_F1_G  ;
and1_14603: n_16148 <=  gnd;
delay_14604: n_16149  <= TRANSPORT clk  ;
filter_14605: FILTER_a8237

    PORT MAP (IN1 => n_16149, Y => a_SCH2BWORDOUT_F1_G_aCLK);
dff_14606: DFF_a8237

    PORT MAP ( D => a_EQ963, CLK => a_SCH1BWORDOUT_F0_G_aCLK, CLRN => a_SCH1BWORDOUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F0_G);
inv_14607: a_SCH1BWORDOUT_F0_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14608: a_EQ963 <=  n_16157  XOR n_16164;
or2_14609: n_16157 <=  n_16158  OR n_16161;
and2_14610: n_16158 <=  n_16159  AND n_16160;
inv_14611: n_16159  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_14612: n_16160  <= TRANSPORT dbin(0)  ;
and2_14613: n_16161 <=  n_16162  AND n_16163;
delay_14614: n_16162  <= TRANSPORT a_N2576_aNOT  ;
delay_14615: n_16163  <= TRANSPORT a_SCH1BWORDOUT_F0_G  ;
and1_14616: n_16164 <=  gnd;
delay_14617: n_16165  <= TRANSPORT clk  ;
filter_14618: FILTER_a8237

    PORT MAP (IN1 => n_16165, Y => a_SCH1BWORDOUT_F0_G_aCLK);
delay_14619: a_N2353  <= TRANSPORT a_EQ557  ;
xor2_14620: a_EQ557 <=  n_16168  XOR n_16177;
or4_14621: n_16168 <=  n_16169  OR n_16171  OR n_16173  OR n_16175;
and1_14622: n_16169 <=  n_16170;
inv_14623: n_16170  <= TRANSPORT NOT ain(0)  ;
and1_14624: n_16171 <=  n_16172;
delay_14625: n_16172  <= TRANSPORT ain(3)  ;
and1_14626: n_16173 <=  n_16174;
delay_14627: n_16174  <= TRANSPORT ain(2)  ;
and1_14628: n_16175 <=  n_16176;
delay_14629: n_16176  <= TRANSPORT ain(1)  ;
and1_14630: n_16177 <=  gnd;
delay_14631: a_N2578_aNOT  <= TRANSPORT a_EQ630  ;
xor2_14632: a_EQ630 <=  n_16179  XOR n_16184;
or2_14633: n_16179 <=  n_16180  OR n_16182;
and1_14634: n_16180 <=  n_16181;
delay_14635: n_16181  <= TRANSPORT a_N2353  ;
and1_14636: n_16182 <=  n_16183;
delay_14637: n_16183  <= TRANSPORT a_LC6_D6  ;
and1_14638: n_16184 <=  gnd;
dff_14639: DFF_a8237

    PORT MAP ( D => a_EQ900, CLK => a_SCH0BWORDOUT_F1_G_aCLK, CLRN => a_SCH0BWORDOUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F1_G);
inv_14640: a_SCH0BWORDOUT_F1_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14641: a_EQ900 <=  n_16191  XOR n_16198;
or2_14642: n_16191 <=  n_16192  OR n_16195;
and2_14643: n_16192 <=  n_16193  AND n_16194;
inv_14644: n_16193  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_14645: n_16194  <= TRANSPORT dbin(1)  ;
and2_14646: n_16195 <=  n_16196  AND n_16197;
delay_14647: n_16196  <= TRANSPORT a_N2578_aNOT  ;
delay_14648: n_16197  <= TRANSPORT a_SCH0BWORDOUT_F1_G  ;
and1_14649: n_16198 <=  gnd;
delay_14650: n_16199  <= TRANSPORT clk  ;
filter_14651: FILTER_a8237

    PORT MAP (IN1 => n_16199, Y => a_SCH0BWORDOUT_F1_G_aCLK);
dff_14652: DFF_a8237

    PORT MAP ( D => a_EQ908, CLK => a_SCH0BWORDOUT_F9_G_aCLK, CLRN => a_SCH0BWORDOUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F9_G);
inv_14653: a_SCH0BWORDOUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14654: a_EQ908 <=  n_16207  XOR n_16218;
or3_14655: n_16207 <=  n_16208  OR n_16212  OR n_16215;
and3_14656: n_16208 <=  n_16209  AND n_16210  AND n_16211;
inv_14657: n_16209  <= TRANSPORT NOT a_LC3_D22  ;
inv_14658: n_16210  <= TRANSPORT NOT a_N2353  ;
delay_14659: n_16211  <= TRANSPORT dbin(1)  ;
and2_14660: n_16212 <=  n_16213  AND n_16214;
delay_14661: n_16213  <= TRANSPORT a_N2353  ;
delay_14662: n_16214  <= TRANSPORT a_SCH0BWORDOUT_F9_G  ;
and2_14663: n_16215 <=  n_16216  AND n_16217;
delay_14664: n_16216  <= TRANSPORT a_LC3_D22  ;
delay_14665: n_16217  <= TRANSPORT a_SCH0BWORDOUT_F9_G  ;
and1_14666: n_16218 <=  gnd;
delay_14667: n_16219  <= TRANSPORT clk  ;
filter_14668: FILTER_a8237

    PORT MAP (IN1 => n_16219, Y => a_SCH0BWORDOUT_F9_G_aCLK);
dff_14669: DFF_a8237

    PORT MAP ( D => a_EQ1036, CLK => a_SCH2BWORDOUT_F9_G_aCLK, CLRN => a_SCH2BWORDOUT_F9_G_aCLRN,
          PRN => vcc, Q => a_SCH2BWORDOUT_F9_G);
inv_14670: a_SCH2BWORDOUT_F9_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14671: a_EQ1036 <=  n_16227  XOR n_16238;
or3_14672: n_16227 <=  n_16228  OR n_16232  OR n_16235;
and3_14673: n_16228 <=  n_16229  AND n_16230  AND n_16231;
inv_14674: n_16229  <= TRANSPORT NOT a_LC3_D22  ;
inv_14675: n_16230  <= TRANSPORT NOT a_N62_aNOT  ;
delay_14676: n_16231  <= TRANSPORT dbin(1)  ;
and2_14677: n_16232 <=  n_16233  AND n_16234;
delay_14678: n_16233  <= TRANSPORT a_N62_aNOT  ;
delay_14679: n_16234  <= TRANSPORT a_SCH2BWORDOUT_F9_G  ;
and2_14680: n_16235 <=  n_16236  AND n_16237;
delay_14681: n_16236  <= TRANSPORT a_LC3_D22  ;
delay_14682: n_16237  <= TRANSPORT a_SCH2BWORDOUT_F9_G  ;
and1_14683: n_16238 <=  gnd;
delay_14684: n_16239  <= TRANSPORT clk  ;
filter_14685: FILTER_a8237

    PORT MAP (IN1 => n_16239, Y => a_SCH2BWORDOUT_F9_G_aCLK);
dff_14686: DFF_a8237

    PORT MAP ( D => a_EQ965, CLK => a_SCH1BWORDOUT_F2_G_aCLK, CLRN => a_SCH1BWORDOUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F2_G);
inv_14687: a_SCH1BWORDOUT_F2_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14688: a_EQ965 <=  n_16247  XOR n_16254;
or2_14689: n_16247 <=  n_16248  OR n_16251;
and2_14690: n_16248 <=  n_16249  AND n_16250;
inv_14691: n_16249  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_14692: n_16250  <= TRANSPORT dbin(2)  ;
and2_14693: n_16251 <=  n_16252  AND n_16253;
delay_14694: n_16252  <= TRANSPORT a_N2576_aNOT  ;
delay_14695: n_16253  <= TRANSPORT a_SCH1BWORDOUT_F2_G  ;
and1_14696: n_16254 <=  gnd;
delay_14697: n_16255  <= TRANSPORT clk  ;
filter_14698: FILTER_a8237

    PORT MAP (IN1 => n_16255, Y => a_SCH1BWORDOUT_F2_G_aCLK);
dff_14699: DFF_a8237

    PORT MAP ( D => a_EQ902, CLK => a_SCH0BWORDOUT_F3_G_aCLK, CLRN => a_SCH0BWORDOUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH0BWORDOUT_F3_G);
inv_14700: a_SCH0BWORDOUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14701: a_EQ902 <=  n_16263  XOR n_16270;
or2_14702: n_16263 <=  n_16264  OR n_16267;
and2_14703: n_16264 <=  n_16265  AND n_16266;
inv_14704: n_16265  <= TRANSPORT NOT a_N2578_aNOT  ;
delay_14705: n_16266  <= TRANSPORT dbin(3)  ;
and2_14706: n_16267 <=  n_16268  AND n_16269;
delay_14707: n_16268  <= TRANSPORT a_N2578_aNOT  ;
delay_14708: n_16269  <= TRANSPORT a_SCH0BWORDOUT_F3_G  ;
and1_14709: n_16270 <=  gnd;
delay_14710: n_16271  <= TRANSPORT clk  ;
filter_14711: FILTER_a8237

    PORT MAP (IN1 => n_16271, Y => a_SCH0BWORDOUT_F3_G_aCLK);
dff_14712: DFF_a8237

    PORT MAP ( D => a_EQ966, CLK => a_SCH1BWORDOUT_F3_G_aCLK, CLRN => a_SCH1BWORDOUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCH1BWORDOUT_F3_G);
inv_14713: a_SCH1BWORDOUT_F3_G_aCLRN  <= TRANSPORT NOT reset  ;
xor2_14714: a_EQ966 <=  n_16279  XOR n_16286;
or2_14715: n_16279 <=  n_16280  OR n_16283;
and2_14716: n_16280 <=  n_16281  AND n_16282;
inv_14717: n_16281  <= TRANSPORT NOT a_N2576_aNOT  ;
delay_14718: n_16282  <= TRANSPORT dbin(3)  ;
and2_14719: n_16283 <=  n_16284  AND n_16285;
delay_14720: n_16284  <= TRANSPORT a_N2576_aNOT  ;
delay_14721: n_16285  <= TRANSPORT a_SCH1BWORDOUT_F3_G  ;
and1_14722: n_16286 <=  gnd;
delay_14723: n_16287  <= TRANSPORT clk  ;
filter_14724: FILTER_a8237

    PORT MAP (IN1 => n_16287, Y => a_SCH1BWORDOUT_F3_G_aCLK);

END Version_1_0;
