// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

module arriagx_hssi_calibration_block (
    clk,
    powerdn,
    enabletestbus,
    calibrationstatus
);

input  clk;
input  powerdn;
input  enabletestbus;
output [4:0] calibrationstatus;

parameter use_continuous_calibration_mode = "false";
parameter rx_calibration_write_test_value = 0;
parameter tx_calibration_write_test_value = 0;
parameter enable_rx_calibration_test_write = "false";
parameter enable_tx_calibration_test_write = "false";
parameter send_rx_calibration_status = "true";

endmodule

