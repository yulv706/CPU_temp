��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc~����B��W�-c8��"���¦|�db�
{��p	{�z�� �`����X'W�=������b�rJqGo���dϮ�L6��@��VEDA�%~
t�S 4�QZ������B�����VM�^�u ���|G0�Wt��b����ԓ��~E!�rjz��
��H�A<[J�E�+�ϊ5v�b��ջ�ANUd? �����ihΕ���}�z�5&n��R�-�c5fɬc��WNL.��*��>�q�����٥ ����"��y6R�(��Q�-��Ɨ�E<.F3��y+ژ�$%I>j��5�IZ� �F�8���$���&} N��4C}�&�'z���ӿ��̓�'Z�MW����S���r2KX�}u����Bu@b�?�ʱ�x�J�B؏�_��R�闚�*YO��<��
��d�E�qe[�[�`9��z�mM��-U�ɓv_�>�p^�e��x����_ 	>��M���5^sũ|d�+����t����a���vmGR�s��U�n�*\�Z!�� U���+n��ڃg??����]���~��[��{��)3a�;�D�ۭMY zt�	x�Xe��!�5���Fz�!�`�(i3_|?k��\�8f���EU���+z�k�����ap!!v*!��sK_���/2=��@��.��L@n��r�iad/�;��Zag??���:�S}^L�u '�����V�Da:������^�%������侖�(+ ���}�!�`�(i3!�`�(i3�g��b�k�H��^���$E�.�T�SQdZ0o�v�����W��4�����)7E�D��,�`��J�~�;�S��(��"]�Z��dZ0o�v��ˎ%Q�Q�z�וy�ˈ�I���y+�L��IŖ��x'L#ׇӭ��!�`�(i3��+�t2�O.$W�qZA��\�${i���~�;w���v.��2�����%�>줧_T���������Fz�!�`�(i3��bW���t7��?��w���i�&9��<��ͻ[$��6��+n��ڃg??���9��xqw$<�L�k��\��7��J��L�͝���_ �KS�)в}��NP�{7��!�`�(i3!�`�(i3{p�y�H�z�SC�%^|/ZT�@���N[�\��|��Oyޕ�����Y�����"��@-+�{��1��ɇ��nC1O*��z�ϧ�����i�Ə���&,��K����p�' ����{��@)v��Uk\��,n����&P��={u�3�j���)E�L"j[�l�r�f��7m�U�$*8����A�����Š΄,�H'u$�~����pC)��L�A��1V�Z5��ܴ>�%�l�}e�P��a�,k�0:S��}1yYZ��� ����@	�1i�myh�~�*�.i,����j�Ə���&,���9�t�' �b!��u�BޘV�� �"2�#Ȱe�!��[OQ�r��W�%-C��om� ��;��dz�'�uIN�/%җ�8����A�׎o�|.�:um �Ļ���p"8M���&[OQ�r��W�%-C��om� ��;�����È�+� �ⴕ���8����A�����;�B0:S��}1PM��!��GS�ɶ�"�����鬕KG�K��5��̻O���)szc_�.�S��'�0����0�4<+��80PS��J�aNSHk&��g�E�H7�81�Ÿr[�c}�sXy�'�H�ׇӭ��!�`�(i3!�`�(i3�p�?�@W{ۧB�qP7m�铲���c3�i_sk.Y.�I�U�:�ƅf���#��+޺' ��nrm؊(�[���~$�B2���m���-��
�8���?�*���\����۠1S-�a��~OҰ�>��?Ԅ��{��+l�utO��7���p✤��6�э����Q{>����D-�����Fz�!�`�(i3!�`�(i3	��j��|��N9����"��wJ�@,����� |ف�'f$�G�#j������:l�h�I1�T�g��� VU��a�Қ��17�i�P�D�K�y؄@�!�`�(i3!�`�(i3.�)�.��� )J�H���"��ʭX�kei�)�%o-�\%��짐�Cq%��k�`�?��<��t!I��G��mO.�w��4܆i��^)7���Y�.���kp!!v*!���O�{�
;����"��ܠSen��I�����˶Q�[�lه�����<�W.��[o�^��Y0R�neײu��ߙ��W�wR�.�c3�i_s/����N4���� �"�R�-�c5f�/�F�A���'=�Ұ�>��?���:�ȋ6�~��c>pRݴ�c"�b2�{������7��U�:�ƅf얔��fG����6���Qz��\{����b2�{������7��U�:�ƅf��o�fy�_���ȃ:#q����De�q/ه�����<�W.��[o�^��dH�M�$/�u��ߙ���¥+_�����|�Enz�<�]iO���<�W.�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN���HR8��ɐ��?u�kظ�����or�}�!�5��Z�T1ۂ�r���x�d��䖯��l����4$��p`Ԡč	g�y���5��gO�q�����f-Q��lKQ1F�o���h�؄)RvYQW�w����|L�P�i.4
�Ǽ
ՍJ��.�W}Opu���A��n����h�99�mv�?�T�u�2�L� il&�<]��b'3��)dj�#@^7&ģM�&yy���S��S�t�o�	ˀ-@�d4̣��[�7�cbp��'#�>-��;�7����?���r��/?�s�m/CO!坭�悬��2a�{:��so�9#T'��nҍ	g�y���5��gO�q�����f-|�bxKҲ��r�D� �m�'4�a��䒟JƓ�����V��늈���+�;�?mP��1U��w�B���`C~>�=�0�u�}�|��Ft
X���?��W��]'��gzL͊�q������W�I��'�+S�hmA��\�v��n蹵��t͌4s+�nye�gW��a;5B5Y+����^B_��+kG��!���Ёy�;ۂ��IÙ=�Hۭ�f"� R���c&;�+�tM6!�'n�^0oL��pN�5����`KE�R�(�Mq{�f��a���Z�.M1�*_��h�V����^ֻ����XP��ȼ�?���$��hP=H�2�+�tM6!�'n�^0o������W�5����`K�={e�jb:JHn��z�����)���%�a��3-���<=�^ֻ����XP��ȵ�d��w����y{¦�W��]'��gzL͊�q��N�p9:O�I��'�t���c���\�v��1�bC/Oy͌4s+�nyA)�[��oZ;5B5Y+�T�����N�+kG���I�	��;ۂ��IÙ=�H�]�h��j/=3\H�.�5�BZUy��\�v��,��M��͌4s+�ny-9"�v8x6q{�f��a�
Ay�9�6>1�*_��h���Q��~��
c�[��0������XP����v<�y�
i˫&3�xy���X�[I��'�<;e�����~��ڹ 	��\�v�Q�����͌4s+�nycfl��6H�r���q�;���'���Xw�j�7��r��&D�:f��:F�X?�g��U-�ea�}�8�4��O��:����ʶ��rHO��c�i��w
��22��X��7�R��	0�W˗0z�cUL_7ݰ�x%y���I�D�[Ø�;�x�Nu�5=��u��ǜ@��^��ץ#�>-��;7ZF����_�V��D��&:n�Z�ɐ��?u�kظ�����or�}�!�5��Z�T1ۂ�r���x�d��䖯��l����4$��p`Ԡč	g�y���5��gO�q�����f-Q��lKQ1F�ħƿ�9c�ew[#K�%�N�����"ڛ������"nz�%�N�����@���,�-��J��F
�PU�\#+��S�M͈�{�P��j.Z��$�sӢ�]3�����c��(rKg!�h��� $��:c+�I���y���OJHn��z���G7���� $����oa��ܛ�	���������IÙ=�H-ߵ'�ѠzM8%�Y~��`�JKݗZ:���'n�^0o����y�]�\�۟�-?�d���&����{ԕ�h7�{`���������������q�z�e�3�ԳN���#t����n{g�P�1[��=��hbV�֎c�q�u�A��o�`Ż�j0��.@.v�:鸸;�����-V��&yy���͵���x���:'�,o�0������]�v�rbp�M>�Z�)˞v}�<�2<@Xȳ�!�3���#^���u��~ \H�}F x>H�|f�-'�(�����Z�,�,utE�խ��;}�[�f�K�+EC���MWU�?
�se�{�z��x� ]
���4]���$`̦�h����0���,�W�B�޹B$~s%��@�:k vl��{�wƄ�{Ƨ\-TX�Rj�+s�!���r�;6��{g�6f.�0�����+�NB�Eo��\�ҋX����@�ڗe'{2e��e0�|��].��'���Xwyd�2�G�Eo��\�ҋX����@�ڗe':�[���Ը|��].��'���Xwyd�2�G�� ��R�%��ҋX����@�ڗe'��k�t�g�|��].��'���Xwyd�2�G�䴙�t�_<��z��}�Q2�+�Y��)$磨'm�rb��S�)37J*u�"��ȝ�]=.-2R��v���Z鎬�����`�;�33�ǳ��֕�i<e\������0ح �x�$X���LqLT@rm�Q4�x#�+/�pr[c�G۶�8.͐Gdb�����o-�\�٬�a�t�^Q�~g{�P�\<��sg=��Y��G���U1�uO����({�t�{/�+����-����R"�]�&���,�v�?Cc0�욁�o_���M*����97�v�ԯ�`�L�i�@�[,E`t�|��].��'���Xwd�n]N�4p���eq�g��U-�e�M-n����Ց2ˁ��{l�f|��rs�i���%��v�u�=wx4���܂a��Z�ñ���3�g��O���U��Z鎬����)��e������	��m��w���Z鎬���������k��'~����TD��ό���.ӛ�D�a���,�\�I��w��,c�A�L'��a9q't��t�W͆���ג�(�K�c]�y���%JXz�����R"�]�&���,�v�?Cc0�욁�o_���M*����97�v�ԯ�`�L�i�G��mO.����9�dMbZ鎬����)��e��+��9�+WZ�TD��ό���.�y}���
L3�б��4@IE�U��@�ڗe'w�d �����9�dMbZ鎬����)��e���S � �h��6�vg;Je'���XwA���0v7���ca�Ԁ�6�vg;Je'���XwA���0v7��m���D���TD��ό���.�h�76AyW��A�04--@��7BB���3�!�M����0oX�{�#���0�b���,��~�rF)���X�3c/��!�~��zrW�@IE�U��@�ڗe'rF)���X�3c/��!���8>� @IE�U��@�ڗe'rF)���X�3c/��!+ ���֤0@IE�U��@�ڗe'rF)���X�3c/��!S}D��'@IE�U��@�ڗe'rF)���X�3c/��!;,�$% @IE�U��@�ڗe'rF)���X�3c/��!������@IE�U��@�ڗe'rF)���X�3c/��!��I�i=�@IE�U��@�ڗe'rF)���X�3c/��!N�Q��*�@IE�U��@�ڗe'rF)���X�3c/��!���W�Q@IE�U��@�ڗe'rF)���X�3c/��!�gzKJƾ@IE�U��@�ڗe'rF)���X�3c/��!��N��d��@IE�U��@�ڗe'rF)���X�3c/��!jZ�\(��@IE�U��@�ڗe'rF)���X�3c/��!��!Ipd�@IE�U��@�ڗe'rF)���X�3c/��!l�W�櫔@IE�U��@�ڗe'rF)���X�3c/��!�(�~;9p�@IE�U��@�ڗe'rF)���X�3c/��!����}��@IE�U����\u��\W���!���		ןS��=L~΄gO�3f��*����f���,�L�Ǉ���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�ֲ!�
\�S�2y3���u�����!:ޏD�.6�+d�ίp��V�����<o�nïi�JHn��z��k"����_<mDrW�B��ɥ����%�a�HL����rm��U}�	KݗZ:���'n�^0oՈ����a�T��r�m��U}�	z� �j���������d&(C�#�7#^�Vn�^ֻ����XP���e����!�?2^�9R��m� ��?�v=��m�/Z%�m�$��Xo��� ��6"�c+Uު.77��`Z"�Ap]-���O
09��O����ƻ��cbp��'�����C��������8��)h+&_���uK��-�������l����Y6 �p"�5_��UX!�`�(i3Q���n�(t4ޚ"k�$��Xo�� �!��Դ��������%.N2������rAq$��c@���N�)�I��'���ưCv�JDn ��a�]�Ψէ@��O��p��Wp�($2��m �A?�=d,�T=�3�������G�����Gߚ�40���Ψ��F<H�-��*p�m~|�֐��6��Eޒ�������S�hӲ������{ϓ,r�r����G����Ћ�l�T���b\�#vX��!�`�(i3���4]�扅��P0р-1 h��p��]�Lrޛ�F���M�����}���ɀ�����f�!A�>�����$��Xo��s��k4�9Q����!�� U��7w|s���rAq$��cn�0���nCth�_ME�v���I�ἃ��<2� �v\m�~e-}����o�$��Xo�c���KB{[���G��!�`�(i3�j>��i6绰�+���]c��3���L=X�� ��-���G�"�|���=�k[��Ћ�l�Ta+PoC~ �!�+�"�,�>E����Ψ��Fp40�zɈ�$��Xo��xq(V!�`�(i3!�`�(i3�j>��i6��ޖl���ݼ�`�|Lݷ����D�zA�U�Y #��U����$	����	���h����*��@|Jy�Y	�R�ʨ��׸=�z'vh?�����$�As��$_�iبK;��(�'i����x�z]�ۇ5����`KhS����2���B���!�"P8{ϓ,r�r�A��m�����6����8�eH�I��'��Z*9�!�`�(i3�j>��i6P�}�~�q��JG<h��3�8�r���d����&byG�O^}��H�և5����`K��W؟���՟�ҨTQm|��3ĭ��Q�q�v��+BY��9���oL�I�)s�#�=�k�f�:�7�C��zC@���XxvlTiy
T�\X�mǓ$�B����u<��S�P��9=�NH�_��Z�I��'���z:��e�!�`�(i3!�`�(i3Q���n�I���3�5�]qE�&:��^���7��k'�w�����9�Vh��z:��e�!�`�(i3�������{ϓ,r�r�x���:����vܴ
�I�����5����`K�`kl�O"!�`�(i3!�`�(i3���4]�<�Z��c�ν��B͡�2��m �A?U-� M�ˊ�a��׻!�`�(i37w|s���rAq$��cE�Ŧ�������Mׇ5����`K4���ϛ�!�+�!�`�(i3���4]㶘p��Kru}��A�"�b���"v��f�;�>)�p���}<��&�Wz�+�@{fT�1�߽K}��׍����}0�st&���\�vūx`��:�,�qo�,ܛ�	��|��	(���zL͊�q���19TH��@���U@���:��F���V!���IÙ=�H�C&�����&� LK�a�Y�!��.�Ҿ�y���O�*���.�gP�����°��b5(��2�p�P���/�K�"A��>� `�_T���j��gf"�	-7��T�Y��}AR�>~qO�P�H���Y�T�\ ��H_5	���Q�$�k\_x���� ��`A����3c/��!\m�U���H��z���8�n��$���fqL���6��o���+�@{fT�U�L�#_���29a���Q�)r��>�fC�a16�o�3��.�`r���)e�k�j��2��xȆ?K�'H�U�q��&��Op�ե[m��5����]�ql��~������ y��!���V�7�	��k��@U8�;5B5Y+� �i7�sp>�.H9���!e����>g��|�����n\�F�9O �?�1���6��V��T�ژ�k��Mf���9���U� ���_j0��.@.���=��s��{`�����#�F���Ig`i�ҋX������S8�	�Ms��3�˷���T�\ ���h�k�����p߷T�!n}y��p�VU��Jm�QA�Q* *e��Q~t ��Ig`i�ҋX����L$�����/'٥��gV�l`�݃�|��].��'���Xw�����C�>�(}%@��7�������{l�f|��:2QYeƈ�=�<�^QP�<�4�8k>6s����]�!��	Ǹ�y85�x3��~�G�
�܍z��T�\ �������>�F����U���>$o?~�d�q�Ƒf����ǳ��>$o?~���C�/7���L>+�@{fT�U�L�#_��H'�t<9�	���K��U�L�#_��f,�GD@�F��qW��Ґ�Yj��2�+~c���<ڧ���3;֍��C�0�i���R��������dL/zV6N4];ˍH�T֟��Bɬ�¦06gM��oP�8���mt��J3؅��FJ��o�C���j0e>r��;�L�|Hj�GD@�F��q*������*lw?��.H9���bP%�uk�؅��FJ��o�C���j��Ǌ�C�����G�Zi-+Q�"�"�=I
Up�]�!��	Ǹ�y85���Vԓ4��[Ø�;�x��Cҷ��e�ˇ�h��<�W�.�P�;DxHB�� "SI���}�]�!��\��'����+7�lI�S�)37J*u�,�JL�����h��R*�&�(��ҋX����L$�����/'٥��gVؤ#�F�#g�]�!���\B��VV�HL�����bQ���'���Xw�����C��FD�(����{l�f|��:2QYeƈ�c�Z�~��w��>'�ҋX����L$�����/�Mv!���xi�ȳ:8Y�]�!���\B��V�W���
�TD���rs�i��ZIp����M�O��6a(􆿳�e�&���6"���
w��(�
t�������2����U�p��
���)��ZbMHmH��R�Q��=z5��*t���S������
�=K1������S���W�5��� ��7��?2^�9Ͱ���*U�&yy�6���:m�ޥ0D�������m�Q���n�UacX�sl\�8䮨�����p�n�ݚ�Н�WK�B�2��5D܅��yu@�Z�&v.��RE�8�(��wC������+q�������Z,'��wO�/ʸ�~{'ia9�j���B�<Vo�eo����ߪ��w|#9����eR���`��c�@+�b5(��2�p�P���/˶����jf׿q�5BO�*����!�2�L: ��ME�$��ҋl9�j���BG+�`'�z�@kSQ����I5��L+lcbp��'�\��I�pD�����y�b5(��2�p�P���/M�UhE�w��E����FO�*����!�2�L:���1��e�"B��$"�s����2��L*P��U@De�0
A���]/�oRA�'�ա	[�*��?l�ϑ��[�ֽ�?!����n	l��)�Z(��/1v.��nq��63�p����nZ8-B:��|}O�*����+BY��9�i_P�@��;U�Qb�|#9���!�`�(i3�E��WC`V��uH��f��WY�;Kcbp��'��ŀk�\e�V
Y>#4q�����f-��9�K�1�r��g},�8���/��+̬was�
���)�b���"v�$�NeG'���E_�OC/률��ͽ�TaN���:YJ�cRC��!�`�(i3)Q*_���x�6�.�)�#�۸7n!�`�(i3j��ԁÆ���ߎ���ղ���<��ᶹ�;d,�ﶉ��eŞ�����j][3�X��ᢒ����u�����!: Kq�ƑYr��ڒ7��ʇ8[�rV@�\��h]���3��Z��(8�q���N:��,��g�7�ː<����}c8sD��+BY��9��!��	=?��FCC3���Øf��x�3#�:[z$��SP��`�.�P{>��ܐ�~w�	s"�֙"W���_K�RP��r\�z��`Ø��NF x>H�|vd����bHl���G�К(�V����p����K�t�1PUaB�s�9)�����m���{�bHl������ڂѦ~;�&}/����K�t�1PUaB�s�9)�����m���{��:: u���� +��X�����Lb!��u�$W��:�m9yI'�t{b@���p��1~��P����9�^�4�9�j���B-�F~>;mn��#�8�D���V4J&)��ٰ���J	��N2v{E�P���^���9$^�����\o�LCd��z��Vի�ٙ�D�s��Uڍ YKf"�	-7���Q�
N =�9��>�������q�}�owђN�~R�wX�������<H�T �����S�	RN&�p�)�3��s�U������6t/�?i�?���5-}�G�1�؇�bu�U�^>��9�j���Byy	}�Y�Aj�X����Е�Ƕ O�YL�P���?i�?���5-}�G��҂r;�1�2h~�wmcbp��'6C��\FTXm2$�mH�Ƨ5l{�dZ0o�v�?�iĉ-�H4!���0b!��u�B���p/.��N*&J%��T���e�F�V��f"�	-7����s�K��g��U-�e�Y%���I�,u9
\_@~�B՟�Ͼ�[�7���DQwF�Q�q�v��+BY��9舩�&t3�$�8���/�К�=M?��v�����h��%a��4�I!s8y5��Ĳ�<����e�F�V��f"�	-7����s�K��g��U-�e�Y%���I�,u9
\_@~�B՟�[��1	�%Դ���l�J�9!�J^�vtiDLq�����f-��9�K�1�ᵉ3���ټ*w2�56b!��u�B���p/.��N*&J��Г�N�;e�a@�}Ř^�vtiDLq�����f-��9�K�1�ᵉ3������^��%fŀ��z���y������qF���	�@�Vw4+��ݩe�F�V��f"�	-7����s�K��g��U-�eן�-�Q�Z%fŀ��z���y������qF���D�ԗ�CW	�h�|����l����4�n���xǊ�"JA�LaP|#9���}�
�?��]���ʣ}��R�0�;"��9�{��O7�4J&)��:1�#��ЭIb�ؐb���`y������GI��"�bK�������\���u���vg!)�='��k=�Z4J&)��:1�#��ЭIb�ؐb���`y���1~��P��=�5Z��a�Rw٥#��� @��������d��9�j���B�<Vo�eoB;Ի�/x�R�wX���p2A�����r��F�����1~��P��=�5Z��a��|F�2�cbp��'Ӡ߳A��A�������=?��FCC3|#9���}�
�?��}a�X�`�e�F�V��f"�	-7��.7��?��uJ�����벩��Y����^��%fŀ��z����	3�� "�q��+BY��9��!��	=?��FCC3|#9���}�
�?�D��T�&D-�^%�ף p�P���/\o�LCd�O7̚����]z8/B[�f"�	-7��_�@6ԕ�8x���:̠�&A���T�\ ���X%��>�o�Q��	�]S3\J��;��9�j���Byy	}�Y��<1(f}ظ�����Bk��~�v9�V}�
�?�,�Z��m	��.�>�Vc����{u�=wx�8���/��F���D��CM��ߪ��Q[R�77��"=�������O�u�9h��xl���fPUaB�s�9)�����m���]�A&�CM��ߪ��Q[R�7b!��u��M���ed�>wȉ�jf"�	-7������C���Hm����v��`y���0���2��f��_¿�����16X�'�����8���/�6C��\FT��Z�-��!�z�د��zNׇ�N0���V�8��R�|�"vQ�q�v��+BY��9舩�&t3�$�8���/���E���T�#�FD�V�����d��9�j���B�<Vo�eoB;Ի�/x�R�wX��\o�LCd��c�7c	��9?���cbp��'6C��\FT��Z�-��� Wݒ%L���m�pз�p���Cb!��u�-)}zyF���y��ϐbU`�(�5a~�cbp��'6C��\FT��Z�-��vT &rd�l�G\o�LCd�t{dU'd̈́���z�e�LQ�q�v��+BY��9舩�&t3�$�8���/���E���T������<~|��9$�^%�ף p�P���/�n�G|���Pc��?@W�m!��ʧɓޒ��s�r�_���:` �b��0�u�}�|�5!��@,%fŀ��z�g�S���We�F�V��f"�	-7��_�@6ԕ�8x���:̠�&A���T�\ ���X%��>�oS��o�0K�5�R��V������\y�~��~/��'e����u*w�A\o�LCd�h����0|�E����F���K�t�1PUaB�s�9)�����m���{�%fŀ��z�s�f� N��Z^+�U�f"�	-7���Q�
N =�u�=wx4���܂��E���T�����@�k�4A݌nNQ�Nw�x�S/Q�ǀ���'t��t�W�$����v�}�
�?�4'�u��vn�J	��r3[W��Pf�K�+EC�M�_�����&���,�v�x�*aE��������H$�DZ� BޘV�� �`�M7Э�=9$Z/�y�eV�PD�$����O�{�������E�z�I�,u9
\_���s,�Uw4J&)��:1�#���,�%kn��'t��t�W�$����v�}�
�?����A��
9���Zf"�	-7���Q�
N =�u�=wx4���܂��E���T��B�.�������L`4J&)��:1�#��ЭIb�ؐb���`y���1~��P��}��\�{��������9�j���B�<Vo�eoB;Ի�/x�R�wX��\o�LCd�sj�D���Z���N`'4J&)��͈H��<����Oo3��$��nt��z8�J�1~��P��\���<�E�l����4�n���xǊPUaB�s�9)�����m���^��K=J��(���B��X�/R�ό���.��������o�x*�+��	ˉ�I-��*��=@r�]3�tx�������*'�M��
'W��){9�h���a�d�٣��c�A�L'̙ch� 5A�
c�[���ߪ��wQR�u9���\o�LCd�c���e�hΤ�`��rs�i��O��#$v'J�B��_Ma�~��MM
��,=�X%��>�o�O��S�wSx�lޞ��rs�i��H���GR�>~qO�P:��`�X�O�g��U-�enJa:�/�m�:��Q?����i�[G=3k�)�� -�`�q���U�1~��P��4a�5>.}V�v�/e�tn���2�u�d�٣��>����C�m�:��Q?����i�[�����0�]�!��"��C����t�����dZ0o�vʂ�M�aQY�{'%sgeߪ�{����Z)��&�t5<�m�1!e�g��U-�eQ[׊}�*���b�,�C�A��-���Ն8X1���}�
�?���s�6/�3�֩l�z4J&)��ٰ���J	D���D��&�y"�
A��~ӬDh�Y�l����4��$����7���ko<��&�Z�^�vtiDL@���p��1~��P��}�|Q�f�1���?���^��k� ʞ���}�
�?�o?Y��ԣ85�"�4J&)��ٰ���J	D���D��F�2�j�����U$?�l����4��$����7���ko<�s�r��7���87�
@���p��1~��P��}�|Q�f���0��[b������� ʞ���}�
�?��bw*�-4������\^�vtiDL@���p��1~��P�晤D����s�r��7׿q�5B�l����4�8l����5�p�?� X֎�<��nM��2��gj�'���Xw��E���T��e<1����rV��%�I�Y {l���z^�j\w��0]}�
�?���e����d{���<�������_��
V���>����C�5-}�G�ZT��r{t�/>�?�K!P��Z鎬��������l�����h�hlf!�����<��nM��2��gj�'���Xw��E���T��#���p�鑙粨[�^.�!�_�� 6ό���.�\o�LCd�h{�4w���B���M�-�^.�!�_�� 6ό���.�\o�LCd��Kz�������R[.C������D@c�qt��q���U����GI��"�㴋�Y��!�`�(i3���^��k�$^�����\o�LCd������Ow����1��g�7�"���ʷ��&T��L��6C��\FT�"������p�)�3����38�v���N,[��?�0vxV7�f�7�~q��
dy�~J��G���;/��O �\o�LCd�%*���a��Pg�U�p�P���/��ٴ��{�G��ͫ������:[2.��y�5��dQ'ד�L5ӥ���-���f����Oo;����+�L��J����^lC��ۺ_~?bD�Y:�
�zq�����Z���%;_."
pQ�d�kGQ��Q�ӃT����3���ߴ�t��X~�+q�2~�'J|��-[�v:v�B�_����\�j��Ȣ��@$˺/t��꫕qŧo��K�O��PJ'�`q�'�]�o Oag��!ģ{v����;��68+J�!��Y�)_��@{�& �^��{5F.ō~EMqş���Oܢ�7�Q4�o�pv(������b�_G�KҨL*�ї�>EtГ��lW̠p�:���U���jt|W����F����2�A����KC����%5�Ψ�FQ�03������<�6ݥ5����e�n�xdɨu �䆡X�dr�jf'��H������V���
���F:_ʣX`��_/��IC:GMG�2�3�A�E'��_�߫&�x�n��ؗ���T��@�#���4t�Ѱ�	/~#�� ��{\o|�����d��lnSJ,����#v�<S�IS�߰A�j�* ��ţ#g;UC����*�������T�)�}�����T��.��W����-���3�� ���kѶ���� lo�kxT:b�*������)�-V���̢�7�1��mbѿ'l���c ���m}�2�y�&�Q+.�����0\�-�^���f�RUw����Q�h�ȓ�iӚ/��Ϥk�;��|B}ø��y�w���H1��@�	��h`����Y-��J��׍���ebCb��Q�-�=p���BC?T�׷eh��S�t_-"iG���9�E�\����8�i�`!31u��dN�)�+'0W��^qXF�����z�1�b$E�D_��Gɋ|5���F��S�?\�ڏ �6n�N�G��|��tG�J����	4T���\�nƨP�ʱ:��Ԩ�\�"ߗtl%�]Y�%���Ádo�d�x��u�5!��g�-��7� 6,�Bf�4��%a<��A���0G3��D��;|Lҹ�s3>zTX�!{��emQʧ�>=B/���d}��[�ƭM��g������Hhqu!���5�Nn���4L"�+�va��2kYD��ʗ��'aOދK-\��$-��Ǡ٥cX@n��%1��ڒTs��w���n��뾦���s��%�u�5d�v[�����fA:z��1f���Ol,=����ꆆmaO��«���c7�S�!��ɑ4Y��u�	"Ocbղ%��������:z(\������ݮ��a�=��d%�Z9 �VL�(\&ݣ(y�ט9��V�9K-W�Ǝ����k�*�.�a�n'�,+$\�M�\ȍ�UD�����Z�קd:�Q^S�^9�
�8kp8MY!K�Y-�¯,��)�Ȭ���g��o��f��̎�4I�_�$�!�[����_�r�e
�x�����ƹ1$.:H�Zͅ��<i&����С)ݲ��R����_�r�eK6��:)9�oR�:S.$.:H�Z�&�'�n�e��i]�j(������_�r�e�m09��C���,�Y�U7k?���d:�Q^S�v|�:�ga�\A�h�
�{Pa�{��+t���P�<d��'R=�>��~�˶�H\�����+t���PF	V	5�rܪ��L���B�NV��	��yX+��o} G��.��rb_6XC���d�k���>���;?d������X.S�����W�����C2+5�"��R�)��<|k�݈�x�������yM��ӡC	^����K��hbV�֎c�W�ƙb�;��5jjM詧0�};�k�Īy�B,�.�*���L$��r�+i�J"$��M���'��.�*���s�r��7�-S�\��t޽{�R_�Ԥ�8!7���8Å��=��h�@;���!���J..�E���?��)(�"�ސE}yޱ;��|B�����,
�x��q%DA<���i���ø�_�r�e|�5��~����M�Y���R����_�r�eK6��:)9�q%DA<����e����d�_�r�e�/��5F����_��������_�r�e�m09��C8MY!K�Y-�¯,��)�Ȭ���+t���Piиs� ���)�d˒{Pa�{��+t���P�<d��'R=���|��%��l�Y�rاd:�Q^S�q۽��h�H���j�r��)���к��B�NV��	��y ��f"�$�!����L�����O�ʬ�'����A��(aMq�P���ט�)Q��b��j��ʹ��`6��Ig�{	#�!�T�.�J��:�������A9\>���|�>G��l*��nm����M���kXb8�BJ�֙I������ܝ��4L"�#VP1M�/rt,?���;�m�����Y-��+�l��ڸ�>fJ�)�,ړ=��Y�Rz�����H��AJ6`{x�fr��[�nR*�Px_/�Z�s�c��L53�����S���=��
g��bL�%s�T3��Jj����E�� e��O/Ԕ��d����Jbަ�N�C����Ыl����%�zC|�L����em���K&ߴ�?ρ�o�&�����b�Dz�A4��rsM�R�Zq����ڒ/�� X�]o��ւ
���uS��K��*�g0���ZùMdA�<��U?�)�}��r
�?�H�G�O� .Ќ��ˣ��Pΐ��W��zN�[(!�N�n�� V��>l+� ���L��ߨ�Vy��Lp�[��hV=������~�b"���$D@P�}��SY1�j�f?C�ms�~�E����	ݔ�������������&Y��V�'��С������$}%��oR��ן�/��-ށ� ��*lxi#�3��|��4-�Q�p����i�7-ڍ�mI�ｘA ��
�A�m�Ìw��$����r�9�>���y��&�/|h&jquP�������L<2<����*�|lC�y�ZDU�.�S�<���壦Zw��!#��]h��eh��c:���6��@Ő��tϓ�g�I�*)�W
:�D1Fp4���Y-��+�l��ڸB��=#�f���{85$_��X�
8�Y�6��_���i:[d�d�6T!a~�$�G�Ep��f�1�v���k�"�$������:�� ���ѡ4\�O	�k��Q\�_q���ռ�R-j"���f���8�cT��T�k��Sf,oN�;�lL�r�?�����+�[i½�0jM�Q��V�N�,�V�RDFR7����;8����Cos�a��!�<���CvU��}��h�I�+������cj1�kD�t�Sj̆��=�f�	�g��ai97���W�H�E\��)����>֐����u�^���i���ø2��gL�b�~����@2�Ʋ��O�	d��:.�{Ѯ�w�,��4ҁ�����~�P��@�f��})&�2{t�/>�?�v�.���u-���[���y�ZDU�.��2��[�rR�Z3�@��t+�6�)����S,f�z�x��F��;�I�8��I��d_���]u-��m�38����̕�Іi��?��^.�!���딃�ϧd:�Q^S�"VP�D��t�=o$J<���u�� ��e��a�������cj1�kD�t�Sj̆��]'���ǰ��x�w{�)e��$�В{��� ����/��$���I�AZ��B�鬽������� M���獨e����d{���<���MwBLLPL5?dK�=o?Y�������✚�s���i���O�	d��_�ݏ���?�W/)G���[�����|\��_w��������x�w{�)e��$�В{��� ����/��$���I�AZА	����Y3�i��� M��������{���<���MwBLLPL5?dK�=o?Y���ܭ\WO|G���O�n��b�O�	d��_�ݏ��2ݍ��B�ɽ,�I�2��/�ΐ��4����wOT�&+D��dv��oTN��'���us⥋:����bU��]�Hqr�02��gL�b�~���Hqr�0{���<���MwBLLPL5?dK�=o?Y����s�t�0���Kcg� �|y
k��e��a�������cj1�kD�������r�y����O��(���9�����m�!�"��:�ޣ���K�ڼ��OY�b�s8�)C�cZe���Վ���a(�鑙粨[�^.�!���딃�ϧd:�Q^S�v|�:�ga�\A�h�
��W<�r�I�Y {l,R�������[����0�%����M ���wOT�&+D��dv��oTN��'���us⥋:����bU��]�0����ڠ�a(��R�� M����>��~�˶.�<���aI�Y {ls�]�y/�(���8�/
�!�[�����C�b����}��A<��nM��nx��V�[��JDD�>RT�>'W���y�l��N�PΚ��_̓ 1B$�sp֟kh�j\s�U&�J�0���rq��Ϙ��c�Y���TO�Rh�|�������5(>��m{���<���MwBLLPL5?dK�=o?Y���9�?s�U/�9�%�����7�t4@�<��nM��N�&5����t�^�1�?�d���&��6,sN��tsb�=��h�@��:zM�M�sm��t�S~V]Ŧ�)�@\��PQń�D����	X%+I�$�l'�7��ܓ��;�4����\���V�I�f���r 	�W��{��.%�8p��,]�U��aq���<�{�!���"����_�wS6j�"Hs�4H�O����u�	"Ocbղ%�zQ0u 7�2�����Vc2�����Vc2�����Vc2�����Vcu���2s?L+�I��nQ�(L	��k
fZpxk['�Y9�GKP�2�����Vc2�����Vc2�����Vc�F��I|c�,�[`�l�������4���c�,�[`�l�����f׿����q�>�Y�V�W|�B�I:׷�F׫�J��l� �[��׍��������֡�\�<7�X�e����]��m�n������"���P�`m��';��?2^�9<o�nïi��n�5�F�^hq��:f��3\z'=юbG�����m�/��}�Nr}|���?I
�x���>T��|b�)_O||�5��~�������۞h�G��׿���4G�ܝ�j�Kӕ3���w%Wze�,���q|��&I��d�q��*�؝��6Q;�im����1��ųcD����mީ29a���QU��nZ��v�5j��i7W�wI>NZ����e��X�e�]y�p���ҟ�
c�[��?�n�x��2�Y��hk�o	���^�w�D��_�\�!�_b�ȟ{�z|j�pn�Y?v�<�7�gI��f:)��1�l�Ui���2��Ȅ&N9Sc)|/k�$55�����z�G��U��G�nԸ��zx�8��6^h&',m�	%�P=ZĚ_���p�ɚ
���;�+p�T�~p�ܩv�0�H5MT!K̡g��b��y?����,\ަ�It*���1����nU��X|Qeu��<̵�U�~Q
�J��B�逫��E��̊�R�@Q��oL젡�q�FƈxN��b�@�����M:��2�;�琾BT��f��2R
�x�Q'��0=V��T<�t�SK��s���1�J���3ճ�i
E���G���N��з���R6�.�3��P�́	P6���˄Y�y�"��N�\:����G���NC'0��<��	6���7�"<��B�q|������U"����I��恔���_Ek��y6���?c����I�7�
?q(f�7S�[��m %��짐ck�[d
4_N*D$H_:t���\�L29:(��������
�SN� :�]4պ��@�����:4�U��[ھ��(=g�O���ݴ�M�h�KX��ik0����$<u]9�#�I�X��WG ��xұs��'�q|̿��ۨs0�f;[���xұs��'�q|�8�8����f;[���xұs��'�q|��q9+t�}ǆQV��Ѩ�f?�R������~��a�Ni���Q���
�x��Y�5��-M�O��~�Ѩ�f?�R��M�X�i��ċ�!-M�O��~��D�$0�Ʀ�|þM���������o�]K`+�0��o)cn
V~$�K�"A���v�/e�1z��y�n��뾦�Xl��]�k��3�%�-��j�L���<cut�}^��Hp9���&�(5�;2i�]�C*3���,��e0H�r���d�゗��Ut�\��0�=�Ҷt��N\®�>�R>��Z�c�Z�~��k��;���:���rU�&"��С�⍇������:��KY�[b%Ɨ��0�=�Ҷt��N\®�>�R>��Z�c�Z�~��k��;���:���rU�&"��С�8���$���:��KY׏�����M��a�z6�T�G�`�]08Ӱn�c�$��#�Y���e z�"VP�D��tKc��8�X��WG ���K�"A���v�/e�#;��v�˼+���8�:䩒=]'�D�$0������t5i��ċ�!-M�O��~��B<�q��V�i@�zP��	���C����i�[G=3k�){���h ���i�[G=3k�)���<���"x(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vx��:+Fwae��%;��I2�����Vc2�����Vc2�����Vc2�����Vc�������(�䏓O(6�l��4�?V6��2el��ԃ��tgF x>H�|x�a1��Ry����ڂ�Į��P��(ewL���G"�֙"W�X�����L��&�p�ڵ�2~�����)�\lIɿ���I)�
�\7Q���(���x�Ms�JW {B�ĜTQ�q�v��+BY��9��!��	"G����d��I�v��Q���(���x�Ms�JNUtԸ���M��)s�K�+EC��f16�LX���S��?�ޭ�;���|�c!L e�~�WcQ����%�sf�|�Ǯ|�O]R`��w���D�0��/3Q�L��lA�ߛ�M�5E�Ŧ���sm|{�!�`�(i3i�y���w������Nn�=z�Cr��jF�����D�i��K�O��S�����u1!�`�(i3F x>H�|��5��yQo�	�N�$"�gy��A��7�Q_�X����h@�ԽVA�ڦ�c4��5'J�Ļ��\IK�yEN�h��M_��֋b��-c#��^	���b�,���shG�����ئ6]o��&7��!�`�(i3
�2�n/f�X�����\f�W6�����D�0��D�fۢB�ɿ���I	�ߏ��F^	�8G[���ˡ��w�:5A��pbp� ,���֥�B^bp� ,���֥�B^��6�p���v��A��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�Z�c/�n�1��i���������LPU9����� S=?l�x���sG���-the�������������@;�!�`�(i3!�`�(i30��w?�h��(Z+�<Vo�eo��l��o���b�`S�|{�]��>�gs�A!�`�(i3!�`�(i3<��Q��\��jT�):1�#���,�%kn�ؼ��J�@-��
<KS�[!�`�(i3!�`�(i3�022��9cbp��'Ӡ߳A��A"�= �魌���QE��!�`�(i3!�`�(i3!�`�(i3F3���%Ff"�	-7���Q�
N =�OƋ.]$j*��|듀�
��Q�# 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�3��V�~�A��j/������8y�Q7TE�ٞ7��A��
,�\��'B�U�s���O.C��|#HK����R�܎/����h7���������l�$><��.pܰ;Ȼs���ݚ�Н�9uC:A�~D����n�
�Ġ����G秸�7�9����M�+�ݕ``kfĉ>99��A0ok����ܐ�}�Y_sĝ���09q6]�ŕ_���sBU��L��?J2��}dy2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl���eh��2B�ಔ��\�M���5^sH�<P��1
�H����KodZ0o�v��&��a
/k�ݻ��q���bY0�,\ަ�It*���1����nU��X|Qeu��<�����v)��&�t5��(���M�o��{~7��%��6�8�}��� �w�Ve���y�j\V�7�	��k��@U8���Gw���;1?�[F�sp֟kh����bU^�����|.��b��F�I5!���Id���N��w�Ve�O9G���0�^�A���P?�Ӧ��Z��zH����I�!3���r=Q�\Ih���X �IF�\� s��x�[e�P�^�)Qn��� מ�c�ql9�P��:���rU�&"��С҂0KA](�@��]�B�*�)FV�i@�zPw�4
Qx.��4��҄E[��
&�>�(}%@��7�����rH��i�׻�v�/e��Y0R�ne�so��%����v�/e��w�WL$�~$�q����!��ZB QR�(�-EW2���|�F�Â�&�V�k;��7O�2�l���T�h���X ��*#�IQ܋i����n�Տ�͖N���y������qF����U�4��BۣV:�v�Ӧ,\ަ�It�XF�P�B�6��t�	e���Fz�!�`�(i3!�`�(i3!�`�(i3k��,�́�$�gZh6�8�\���h��%a-K����B���_��P!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3v��+���Q:Z.�M�L$��r�+Q����:KG!�`�(i3!�`�(i3!�`�(i3!�`�(i3�͈&�15I��Bb�z -)}zyF���y��ϐbU�"�O��!�`�(i3!�`�(i3!�`�(i3!�`�(i3G����?>�SC�?�$09q6]�M@C�h���]ȷ���(_o�dZ ���y������qF���J��*`�X�~u�j�@~�B՟�[��1	�%Դ���B��+��!cft
�**�����<˫{�
Zv4=��/!�`�(i3!�`�(i3!�`�(i3�_��������<F�T�Q_o�dZ ���y������qF���ô���2xDp��T�)�k1+!�`�(i3!�`�(i3!�`�(i3!�`�(i3���#{Eb�M�r�kZ�g��o�=�Ž�Ӡ!ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����+E:Sy�Kt��SہS=�:B�cC)yׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3"1��y����Q��4gAkT�s�O��-�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g��B�~l�X;p`�B���p/.��N*&J6rT�Xk:)���2�CK2��@:�s	�i�K����������ը�k:)���2�h�AR��j�QIkAI��������`k�@���t!�`�(i3!�`�(i3!�`�(i3,\ͨ܉p����O,8�?�и���]���ʣ}��X�=1����xDp��T�)�k1+!�`�(i3!�`�(i3!�`�(i3!�`�(i3���#{Eb�M�r�kZ�g��o�=�Ž�Ӡ!ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�����+E:Sy�Kt��SہS=�:B�cC)yׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3"1��y����Q��4gAkT�s�O��-�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g��B�~l�X;p`�B���p/.��N*&J��Г�N�;l�J�9!�Jv��؄aX�B���p/.��N*&J�3�������G������<6��<
f~$ :�Q;�im������3KT!�`�(i3!�`�(i3!�`�(i3�q�9�ͭ���t��˳m�)^�w�_y�AN��K������Np������$#z�*�fH*/�<sȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3$�H���s.�vL<���zj�������1��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3C����|����2�2&O��4�q^�5�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3Zd�N��V:琉��{�U�����sȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3�!��(Ot��5�NP��\���u�;r�6�&{�`��Ҝ~�.״�8�FI�g�M���y������qF���%���C�ۅ� o������S���ƃ�8ׇӭ��!�`�(i3!�`�(i3!�`�(i3��+qсH���0���d�Pq�@~�B՟D��Wp������H����Fz�!�`�(i3!�`�(i3!�`�(i3!�`�(i3����0�X�)Î��C<��10�i}�eS�zTg�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3<9�i�|��}jz�R�ޤ-�N~�]�{�@T���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3>��P���t�ɴ���&�a,�񟃧���Fz�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�O���/�6�8�\���h��%ad�nu�U���й�lK����a�R����6���*����Y�����~��n��� 00�7��W`�n|s�)>cv��k���.a1�&��-�hR�5y ���|4�)?0Qp�&�%)!i~O.C�ׇӭ�ыe�䭫��;���cS�)��&�t5p��HM�e��Cҷ��e��)G�J�cbp��'@
9��y������1�R��Kl���b\�#��	�p2�]�<�!�`�(i3�]���ʣ}���	�a�a�bP�)R��hSׇӭ��btg��|�@~�B՟�Ͼ�[�7�}� ��5S�D�0V���%>�rG�u�ݶd�;�jmT�#E��'�}���ɀ�&�&�IE��"X��[m��I-��]��TM���K�+EC�'=�\��6rT�Xk:)���2��R��Kl���b\�#��	�p2�]�<�!�`�(i3�]���ʣ}��r{����JDn ��a�;�V�u�AE6����	��x��]���ʣ}��r{����JDn ��a�;�V�u�P��^5HN��R��#�mo����Zj���
���fD�"���b\�#�y�Ya�I��g��U-�e�&|Q{� �\��jT�):1�#���حg�̰����J�~�;�,�oQ6s�IG"\�A��7���s����Pi�#��R����L`���h��%a�p3�d�&H}���uy|����]~�|���T՝� s�#�]jc���Rw٥#���ưCv�JDn ��a�;�V�u�P��^5HN��R��#�mo����Zj���
���fD�"���b\�#�y�Ya�I��g��U-�e�&|Q{� �\��jT�):1�#��Б|2ҟ�,tTXP�e�gh:�:g��ngFW&�`�w�Ve��e5ngY�^3ZiY!�`�(i3B���p/.��N*&J�3�������G����������;��AE6����	��x��]���ʣ}��R�0�;"��9�{���#,؉'��z��fĉ>99����y�"��H����f0���Nf�3k1x��T�/R�-�Aa(􆿳�:pP�l?`�'��P��+BY��9�̑PY��ESC���X�?�"��)��&�t5nU>���gSz�����	iV\bւ�@~�B՟D��Wp�����9U�%�]D8|������#ҽ���;��� d��\���u���vg!)�����T;y�'��z��fĉ>99����y�"��Fr��ja�U�ے
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl���eh��2B�.K���o�)��T_��h����j�n�a����#�q�
DgEou�R��Yy��$ŧ�]"Jׅ��E 
]	6������k����*���sSr�K?K�- ������q��>��h���qK��������@�.x���o!�`�(i3,\ͨ܉p����O,8E�{w�%��짐5��{��#�`H`��t&h�C��!�`�(i3!�`�(i3!�`�(i30X�C1n����s�6/�M�b�J!�`�(i3!�`�(i3!�`�(i3B�`c�}%������R�t�anb@����I�d��ݚ�Н�!�`�(i3!�`�(i3����,֘u��s��V�i@�zP���_�f�?ǉ�=!�`�(i3!�`�(i3�O���/�B!�R.e�>��z&u�'Ʒ���%����UC:�<c�C��v=�����+l��?�P�4�=�*��������!\�'��p��^�zL�,�%��짐5��{��#�`H`���O����O.C�ׇӭ�ѣt4�K��U`y�.N�d{Ĕf>�u�^3ZiY!�`�(i36pG����_�f����4
��R�1�etat�r����>?8�;;���Fz��*�RoZ*q����T;y�'��z��fĉ>99����y�"��Fr��ja�U�ے
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl���eh��2B��kY~,֨��跤="(���a��}���ǉ�Y��8�X��ݚ�3��(�<�����iӒs �CY';��7�ޤ-�N~�]>tƤˌe4��A��
�R�	������� ���!\�'��X���k?�}e�6BCq�.^Pi�#��Ry	i[��I%K6��:)9��B��[�^�����&�Z�5'��|��Vu��r��y	i[��I%
�x���B��[�^�����ӛ��5'��|��V��C�ˤk����l��m��j��~�����\��F���P7�kq�
DgEou�R��Y>�$�F�_'0����ڠu���'ln�m09��C!����H����l�R�p	��fM���^a�4�21�2t��y�eu�j�~�sgѼ���5�����Q���jV�w(}v�qz�}��SہS=Ѧ��hN캧xӍ.��v�/e��Y0R�ne�u]�MP�<�2#��2��v�9��fĉ>99��A0ok��$f��_Ub�$Q���ܛ2߸��S�Ȍ_�,|jԤ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�3��V�~{�����P�ք�ώ�Q��`:���d��	��I�~|��9$]����";`y�.N�d��;e��J_%4\��`l���L�[(�.D�7��Ł\x�"l��F��':`~|��9$]����";`y�.N�d��;e��J_-)}zyF���y��ϐbU���=����<��(�@|�|����!�`�(i3�������l�*#�IQ܋.�S�nL4Gô���2xDp��T����!+�*��A9`"�
��R�1�e�����ը�k:)���2��=���~E��T����B��+��!cft
�**�����<˫{�
Z&�2����!�`�(i3,\ͨ܉p����O,8E�{w�%��짐5��{��#6rT�Xk:)���2�}��o���!�`�(i3!�`�(i3!�`�(i3`�.�M)3YG���Y&�y"�
A�����!�`�(i3!�`�(i3!�`�(i3<9�i�|���E&����K���wS�f�?ǉ�=!�`�(i3!�`�(i3!�`�(i3#�*�5R��a��fv����QX�`!�`�(i3!�`�(i3!�`�(i3�O���/ѧ�i�6cl�J�9!�J�j"Xt�F!�`�(i3!�`�(i3���aR�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl���eh��2B��(�@3l�H���� 7E��^�y����F�-��M�(�d+�'�����_��t��W�+�!��]���I��N���7�¥���Wt��w9ֱ���=鏳��8d�,�Z��m�7Q6�1F�;��?�;��?��������r\�z�_9��o�R�rcJ]�0��0p2��.�=ۡA�qjwu�Z��K�zb�p����	3�q����.q��r�������L0.�L29:(u��v�<fD��%��Q�9�=����.̪����Xz1{��9����W�W,R�����N�(BqO�s�I��f�RM@	C�	-s�*w�!�`�(i3!�`�(i3v���u����~�R)�rޏ���[d��]&s�|��������a�<B� ����M�Yag����g��BK�9������mo1��z�׀�!�`�(i3!�`�(i3��b��\s�$W��:�m9��$#z�*�
��A0���l��cx5����yy�s3�qԿ�!�`�(i3&�XS��n8|C��t��A��
fhQs,�����(�
��R�1�e�Np������$#z�*��2��\% ႅ�a�mI$��
�O.C��|#HK��^�+oI|���� ��1|F x>H�|h:�:g����f���k:)���2�<���H��d�%��l�J�9!�J�@�QV�`�^`H��%�S�<A¡f��� ��1|F x>H�|h:�:g����f���k:)���2����ў�L-M�O��~�,9]�y�b�dZ0o�v��O�z��,�7D�EI{��^D�����d�tð��T�ݚ�Н�ӯ_/T�ŧ�Xz1{��9����W�W,R�����fD�"g����P�Sb"�3k1x��Tl\�m*k�N��0����b\�#��	�p6 -�&���r����	iV\bւ���k�A�����t_!0xm�N�f0���Nf�p<kd�$ʣ'R񔫇9��)�c�D&������A�<q1���~	iV\bւ���k�A��� ��JJ��T��Ě���P��U@Dφ��<�6���?�B�b�4���Na�CLap=��[�O�%���?�
;<���xL<���xB2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������ʐ�;BT�iW����n�G|���Pc��?@W�m!��ʧ��9-�b51��3�������`�$���-�L}WqA	��ı%z=( �m�OQ�£\D�CT;�h���C�b�&����-%4\��`l���"#RW���t���][Te�u�>L�$rK|���џ����h,��_��h�AR��j�QIkAI�������φ������~Wv�|9�!�`�(i3,\ͨ܉p�u�B�bϼ�X;p`�h:�&�f�!�`�(i3!�`�(i3!�`�(i30X�C1n����s�6/�M�b�J!�`�(i3!�`�(i3�)�0��qvZ�`茟D<_��`o�o�ݚ�Н�!�`�(i3!�`�(i3Zd�N��V:琉��{��dE�J��!�`�(i3!�`�(i3�g��B�~l�X;p`����L�Bs�������<;>w�K���s�?�oC:�<c�C��v=���8��H��R������ �l�J7f��]#�g�4�ɨ�A�,�v_ ��K^y���M�-
�k7�+k�t�m��-s�?̏���m�1����}�ю�A��
fhQs,�Mt8w���E]c�%��=Fh�z������Ȇ/[=l%��x$q�ᙠ&�(��!k2�-�*��o(����<mF����>)�>0�")�g�d�ԫ[=�.n�5�����}YBG>��d������MM
��,=*A&-�Ri!�`�(i3RB*�5}��`kl�O"�B� �b��!�`�(i3	iV\bւ�;8n)ͅ��kq�)-�o?Y���b�_A�z!�`�(i3�����!�`�(i3	iV\bւ�m}�F%iJ!��g۹��9�P�[�h�=���]����y��F�Z��8�M_��+3�Љ!�`�(i3���F��O��ݚ�Н���iO�_�FR�f�
%��v��!�`�(i3�?�JY�)�q��ڍ��jVѭ@����l���e
p����ϸ��]��TM���K�+EC��j�Y��r�&T��L��O>������ݚ�Н���iO�_�FR�f�
n��뾦�!�`�(i3��tM��� !�`�(i3�({�+�y��;���b+}y[
�:qEp�;�P�t�5!�`�(i3�EK ��yӧ(BqO�s�8���/�����W�~j��ßn!�b��v��]&��:0!���F��O�i ���=��4����RŚ���>�LKo���x�2 ��4�ve(��yNR��ڮ����A������B�M�5�Ta!;
=Ի��2�f#c~KZ��}/Üy�a
�:v���Z��#g�k������Hh���gY�Ix��Wǖg3ȓ8���/���D�1�#��KO�7`r�}a�X�`���
�C��"X��[R<�0/60H�/8^b��w;��|B�ڮ{�6,�DRM(�e���dH�L�
�D�3dQ;��|B"�J��Ǭ_5)�D����sͧ����P�$�7����,�ǰ0�:��iy�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc1 T�V	��0?|�Pc��?@W�m!��ʧɓޒ��s�r�:�E�\����jXaP��ɂ" �O��W��|�>b\���5������j'.T�n|s�)>+l�utO��#9j�*�AR������[k�#�r��q��SScxo�ߪQ��fV$vHSmH��T�٥��T?,>�y��6�m���c��?��d�����{���R�$c:���y�e���HO��4��d�S`��o�ݥ&N��JDn ��a\��猘�`y�.N�d؝NF�a����  J�X�=1����xDp��T�;V4�E��\d=��¾ȼf���Ն˚�\��6u�=wx����ZqJ*A&-�Ri	iV\bւ���Kf�g73Q��*�q�
DgEou�R��Y��4��҄F���Z�Y�I�_�(������H�LxDp��T��-tN�a�U�/��b�����$h�I$�-��q�\�Y���I�ºg��BK�9�-ײ��IF�\� s��=�����F�fyևM���5^s�.V���x���g��o��8���H���~����W0�]��x@����ܐ�}ć����akQ��fV$vHSmH��T�٥��T]�G���Ƹa�������pU�+��u��Nl�J�9!�J�����E*��,
�;4'�u��v��
�+�Ϻd=��¾ȼ;�jmT�#�]ْ/:�;̲@�.�X8�{H�RtV�^�����+]��¬j� 't��t�W��2U�5;����Yk��	iV\bւ��s+Α�9sD��αt�4Ⱥ�o�g��U-�e�,���6+�fĉ>99��R�V�"�0ɉRa])n#���r������DQ��&�sх;���4A݌nNQ��}Dq�f��5ߧE4��W?�;��!2�͞nOY��a�R�Q�z�וy�C.�����f�aolm�K���p�gI��1�W�^}su�V��M���,�5)��'K�]��¬j� 't��t�W�)����]�5�O�%E#P\�
�=ĭ,���P)��=��h���qK�����������/��f{�ʬ�缆v6�o<5�!�`�(i3!�`�(i3k��,���#Lk�j�~�A*����X��!�`�(i3!�`�(i3!�`�(i3`�.�M)3QDTy�V��P[�$F��|ʏ�ߖ4!�`�(i3!�`�(i3!�`�(i3`�.�M)3QDTy�V���ӛ��f�?ǉ�=!�`�(i3!�`�(i3!�`�(i3�o��Bl�FO-Z�'��Fے�K�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3>��P���t�ɴ���&�a,�񟃧!�`�(i3!�`�(i3!�`�(i3!�`�(i3�;MR&�l���2��i ���=��?�d���&���4h)qe��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hAj�X����DV��0� �l������|�W��	]�	�>[ŷj7�hr����ޓ�x�&bm���ӿ�G��!UL����0Fo�!�M�����i˭�����!\�'��p��@�.g�L
q�
DgEou�R��Y-�*��o(����<ms�� ���L���m�pҥ�՘�'7I/��\]� h�ҩ�Ϭ�F-���(��P0\.���B��rL�`y6��j�2��	��x�4'�u��vn�J	��r��x� �p�my$�N��o�/���;fĉ>99��A0ok����ܐ�}ć����ak9D���o��Mt.K8��2����_��Jh��MkE��p��-�~_�m�À�p��xq���̀���<��@��v{�GvWދ�qc:�rcJ]�0ݫ���Uh1�;��|B���r����_Z�����h�AR��j�QIkAI��������^ �7�}3�d"T��O$>�����w�!�`�(i3���f�MhhjXmRQ���7_]�4"m��1�M]�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�F��*6�&�y"�
A�����!�`�(i3!�`�(i3!�`�(i3HK(�M��43� uZ�x	�����l]�7߈
1���.D�7���&_rm����!�`�(i3!�`�(i3!�`�(i3G����?>�SC�?�$09q6]�� ����/!�`�(i3!�`�(i3!�`�(i3�/��d�$��Eeu��S�V��!X�x1�"�h<9aV��	��y��@$p�m����x���H`�)}�=2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcwz��
��:i^��������_ŭ��@�0f �pC��)Va.��2~�����h�j�t�!+}ԓ傑��ئ6�)�U 
4�('ro��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcwz��
��:i^�������A��
��;e��J_�ǁ�����IR��IF�\� s��ђ*Z����RVM��%��$� )�a����KM��-�t��N\®Z��@�+��U����if��O'�������~�d�'���T�$���z����o8��OƋ.]$��CW	�h�}M,�d�JDn ��a�6�	G_[Z�T�0Zg��BK�9
�fa+^F�ኟ��L�l��� ��1|F x>H�|h:�:g����f���k:)���2�ه� �4�<���|��@�,s�K�
�� o������S���
�C�1h��V�Ҝ�R!�`�(i3!�`�(i3�dv��oTN^q�e7����m���Y7����&���,�v��0�^��ݚ�Н�!�`�(i3!�`�(i3jJ��I��n��i�a�
�x�5��h��!�`�(i3!�`�(i3�͈&�15I��Bb�z IF�\� s�ʸT2p�!�`�(i3!�`�(i3!�`�(i3���(R��E~�Śg�W2���|�Ff�?ǉ�=!�`�(i3!�`�(i3�6zq��J_o�dZ R�$c:���4p���eq�g��U-�ed�$�IF�\� s��t�j��1
f~$ :�Q;�im��5��83�!�`�(i3!�`�(i3�dv��oTN^q�e7����m���b3QyP�h�ݚ�Н�!�`�(i3!�`�(i3���#{Eb�M�r�kZ�����~�r���!�`�(i3!�`�(i3!�`�(i3���)������m���.� f�T����8��*!�`�(i3!�`�(i3!�`�(i3>��P���tw�'�{�{!�`�(i3��_�����}p���V`��!�`�(i3!�`�(i3!�`�(i3]-������FO-ZƐ�%�`�t�q�&V�������n|s�)>+l�utO��#9j�*�A���R�&�۝-/�U�3cה����7���o�m�nRQ&���*���]q�����_��s�֙7�}�!�����A��
�[,J,�R#�� +6qd�N�Luy������`���pF_�<�K��2�O&�zH���u@�W(FOHZ�.�g3Zv���� �ct������~���hc��eV-����1~ҟ���P��Z��m����&���*��µ��da�_��s�֙7�}�!���J���7�����2�=Fh�z����D6�saQ��*��i�벩��Y�O�����X���/��>�.5o�fa���{���w؂��\9�o��R��p
���[�����(����<m�Zj���
�Z�B�ӿ$r)˸�h��(Z+�<Vo�eo�NL�l'*/Üy�a
�N���9��F��|��ujD^k�uQU�.P	HȆH�RtV�^	iV\bւ��$_�[o8[�%��ؿ8���NM���՝� s�#��������A��
�[,J,�R#%��v��!�`�(i3���F��O��;b�-�2�$�)�vx�]��<Jf`��!\�'��$��f :f1 �]C>��ӚH�RtV�^�����+[V��M*�&T��L��[��(��!�`�(i3�t�ho���[=��s����~j^�q�����f-D2�����?�=��)�*����^��!�`�(i3	iV\bւ�~��Mب�'���irU���|e"
�:qEp���e$F�pF_�<�#�jM=)P<�ܓ�Y!�`�(i3$f��_Ub�F�S�1 �HN��R��Gu�"�0�HN��R��4����i ���=��?�d���&�۔%��)���m���]T��hV;�����*�)|/P2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����䎕��4"I��A5��b�>pRݴ�c"1��_���6�o8:4�IF�\� s�]��s�Z�f%$e��?%4\��`l��]��*�x6BCq�.^H�RtV�^��� �l�J�9!�J/�\V,��K��"h��:���rU&X�/(ӠyU�.P	HȆH�RtV�^!+}ԓ� ���췭't��t�W���[�4�f,�rL�`y6�RUAY�"'t��t�W�'�[�®�՝� s�#f���u�[+l=e��0�U+�qbp@����%>�rGO�D mWN�׹���U�_��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9z6����T ����F��|��u���Č��f�R�5�Y�IX0F�M�9�'
�n6BCq�.^H�RtV�^ Fah
8�xm�N�f0���Nf�p<kd�$ʣ'R񔫇9��)�R�
9����^2y9���ݚ�Н��}�W���Hc�[N	K״$(�>g��Ra])n#D�
 D�Hc�[N	K)P<�ܓ�Yfĉ>99��A0ok����ܐ�}ķ�����q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc1 T�V	I"� ����s]bi~�U9�����"n�E��~��Z2��z�fU�^�����Ϩ�V<��1Y~��`�J��xG�"Dd&(C�#�7#^�Vn�k�O�>!�`�(i3!�`�(i3�q�9�ͭ���t��˳Ie���0�D�ػ��DIY�5����Ң��U�t�!�`�(i3!�`�(i3!�`�(i3!�`�(i3p9f~ݬ�n��i�a�
�x�5��h��!�`�(i3!�`�(i3!�`�(i3��>Ո�9�=�8�_y�����H��>�B7Ԅ��!�`�(i3!�`�(i3!�`�(i3
QDD0[���^@R�C<�2#��2B7Ԅ��!�`�(i3!�`�(i3!�`�(i3q�8f�t�tu�$��-v7�"<��B�q|�#�y�
F�S!�`�(i3!�`�(i3!�`�(i3!�`�(i3flY��,��Na�z�N�k��!(=-[Te�u�>L�$rK|�@��]�C���9���V�i@�zPw�4
Qx.f�?ǉ�=!�`�(i3!�`�(i3!�`�(i3JZ��2:��X;p`��+t���P�|!�}۩P!�`�(i3!�`�(i3!�`�(i3�eR�ﬂ\�H
<��is���'�2���B� �2Y)Z:2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�pv��[�\�k�D�\�w0Nj�C�T8n)d�K�ծ?�*h�Jﮨ��������i
f��/�gm�t.�6�o8:4������~����I{r��èV�Zj���
�����~��a�Ni��y;
�R�&�y"�
A�a��Dx�Q��-��������l��w'r����5�����Qx{^4��*m!�`�(i3�/�L�s�jJ�ϋ��-`ƾ��/��5FR]�[�ܒ	��x��ݚ�Н�4����$؃��yi7��SN��,k��e(����;�P�t�5fĉ>99��A0ok����ܐ�}ķ�����q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcwz��
��:i^����or��ݔ�����G�$W��:�m9�@�N���153p��z�:j� ������fH�SrPc��?@W�>C��p!�ss�������k����*���sSr�K?w3�_�]!�`�(i3!�`�(i3�����q�,]���	/�g���̹��
��R�1�e1�؇�bu���!+ٶ��6'�V���R�8@]fy1�@�>{2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������Ak����������+��7�g��Q�;��֞��� �����9qK��[ ����I��!\�'��p��^�zL�,����A��
L�j�=2pөm�@�[@r�/dI$��l�Ig?|յ[+8�hV�6�����:^)��4m>�B�t�c�ѧ���O˿+<b�3&���M[��ޜ�}Dq�f�f�vWb�P't��t�W���[�4�f,�rL�`y6�RUAY�"'t��t�W͢^��/�� c�j�Q�cO�ӽY�'e������:��_i ���=��4�����i_7�P{P��˲��Z�
�x��.���HI��]S�%��èV�Zj���
�_m��<<���H��O잢+`|"l L�BV�����v�ـщ�l�Pp��s�g��Iw8�}�����>�EWz��ُ�&+Ä4����$؃�feV���'�^�����;b�-�2��6h��07o
�x���B��[�^�����ӛ��!��}���џ0S��ϐTZ�1{~�Xy���9����eu�j�~���;��*�5�����Q;Ȼs���ݚ�Н��H������r���܇q|̮���+c�g�d�H�RtV�^!�`�(i3������Hj"X�U��y��)�r��:5A��p
�:qEp'{w#/ B!�`�(i3�	z�5��R�qE?9�,�'��P��+BY��9�`>	�S(c��5%�Jm�#������Y�8HV�,C���Wk���1"��5��K?T��}Dq�f�!�`�(i3�šB)�/�H�,3)��Q�o�8�l^������|e"!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN
�:qEp�;�P�t�5fĉ>99��A0ok����ܐ�}ć����akԱ��+��i���%Ὠ�p���\���`�+N��@O��BK-W�Ǝ����k�*�.�a�n'�,+$\�M�e2܂A1%�#g�k��rV"�I?������m��1"��qG�aYݍ�?�d���&�Ա��+��i���%Ὠ�p���\���`�+N�Y��~:=�Kv��f�F�G���6���U6!w���W�����C�1ȉ��������k�*�.�a�n'�,+$\�M�ӳ�?RZ?=|q��M���rU���6�h3��bӖ������μ�O�nV��	��y����}���H@�{�'IK�L�����d�kⲩ�Αo��p2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�m��O�{��<|��7�"����j��I��+���N���6����e���s�6/��)�}焓>-2H��.�-:��y���I9B,#A������������:i^�����4�r�ӭ�q��JU[��P��'���ǂYJ3Eo?Y����)�}焓&��lm���͎)@�Nk��+t���P&;7�l�\9;Gt���m�_�6ʳGV���i�[G=3k�)�mQ���Mf�^n,N��M&nȹcJ��+�A�wv��؄aX��P�h~T�5�'������SQ�5	@<ӵ?���gY$���H�rg :%ri�$���.Mf�^n,N��M&nȹco?Y��ԧx���i�9Wrb�B�epƽ���+t���P8�=��j>KH�v���"�Uђ2o?Y��Է'�����ƛb�;�Dc�J�L�`�;@��!�EUttl9���R�<lͬ۞h�G����n>���(=g�O�?�C<xWY�K��e�Igg^�`Â��M�Ƿ�>�wN��UDz�w�'�SS������{�T���v��LE�����[�i�R�<lͬ۞h�G��!g�U�g"`z$��S��?�C<xWY�K��e�Igg�R�@�3�0���m����	'����'�SS���L-�yC³ˬy����O�@���E.�R�<lͬ۞h�G�x!2�͝4"|�$�T�?�C<xWY�K��e�Igg�{��E0��C�	7��/�4e�{rF)���X�3c/��!���7�&Nк�h���ޚ�R�<lͬ۞h�G������W�1���4��*{+;����'�SS��F�Y�H�n�n����{
�,m��WPrF)���X�3c/��!��Iq=+I�8�ؕ�+?�R�<lͬ۞h�G�D<��\�zf*�b
�@�L�(�rY��'�SS��/ل�� n����{
Gh;ʹ�[�rF)���X�3c/��!� Rƙ7!���Ɋ�?�C<xWY�K��e�IggTQ�w�m�#�=��E��luVU�簦~09h�i��½G�c'.�h��%��Xcbp��'����Q4KҲ��r�D� �m�'�t�חEʭ�3�Jl�9���v�/���m���B̑!<�!$�Uuy�R�
/��a2&P��6m05YT"F����q��1�:/��8a�B���k�t����]�BƠ���VӴD�(�T�Ù����׉󾶓�^�.�8�7a	��������W;5B5Y+� �i7�sp>����S �=�[T�)���}0�st&���\�vūx`��:�r�^K������О.|��	(���zL͊�q���@F�4��d��X���n5T�n6M�_3#ڸ�l����4�:�����v�~�����9�j���B��S9��c�,�[`����9�dMb�l����4�n���xǊ������ Z�U��c-����"�t���~���b]�iz�9�[vĄ4Ȃ��3Y��Zo���#}|��XH�����,>$<�խ5�PK��e�Igg�1j0���ƸWw�8��pzl��a�o��%H��9�j���B�<Vo�eog���gB��Iz#1�<Td��"X��[�|���M��{_8�Y��=�}�Vݨa'�<� \����K�ek���o�7��K�+EC���>v��T�\ �����^$���w�+��"�A�#���C��iF�(j����OR�JO���Wx�B���6��c"U�_�Z'���s��d�\��MN����!I/�������A��X�@�5��6�l��sХ+�:R 8*�A��jeN�V�����׷eh��S��L�u�RmHX����20)�_h��r��a)�m�d�so�}a�C�ub;�;�����w�?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��Le��	I���]�HЦ��EMW!���4m~�����c-�z��~��D:ǯ3�4���X�E��	�'�J���U�2Gޣסe� <���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+�S�AZL�0hs�A_	�K�o[��mU;լ^<���X�E��>��}z��T��U�oLF�����8�Ɛ�a�����|�Y,�ΊB>���<���Hn
V~$�
�p\,%�0�OvԳ�3뮋ǕB\x;8����l/ǋq܃NQq�cl�j��c��}d�<�Rc$I��h\�7�.�s��a�a���v0�����c���0�K���
�p\,%��b�I.�Ha�
�p\,%��6mN|�?&)�5#�ܸT�~�������� 288���������:�ͽP�$�����Oam�.�H��`�M�ͦ�J {�ú�8�$�N\��
�M����?6�<�U��x]�iQ�V��Ue����{��� >ؓ���zռ5���m�-�M��k�R��9�rn�VpaUv��h�Q�L�6�֠�+�v.V��T��#�-�p�������?�r�J�2E-�Rxp���[0��]8��t 7ڇ\ze���!
��=�*��3P� 288���ȓ���w�SWb$$b�)�oW<���>��Z{��3�����Q�r�yK�9��7�_���.":�!�`�(i3RN�]�5'�b1]�Q:~n�s~��20�OU�TG�eIw{��lD�!�=e�ȩx��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����k��J�Z���>H��L�}�Lqo��L�h� ���ڤU=�v�)�BҺ�)�|�$G^�2u*0��Y�b����{�C!�`�(i3!�`�(i3��Y�H~ XL@3~�����Q_K�WL��<z2��������Wq�`AShV���.�����_q���"�7&!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{q��#�i+����Ó�d+st�I6ȵ��$6�*�yȩ�,���8��	͂'�)�����jryX2�u!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��~��ɳ�GV��)�m�c+
�i��"����vg��i�C$Ԯx�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3rz��G�;����A=&�������3�����Q��ʋ�И_�֠�+��v���V�i�#�-�p��4�= w
��D+���4Y!�`�(i3!�`�(i3!�`�(i3�g/t��5�Y�n!�ƪ�7�t/s�+� 288���� �Z���Wb$$b�)��ˢYۋ!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3RN�]�5'�b1]�Q:~n�s~��20�OU�۾�\��lD�!�Q��S���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����k��J�Z���>H��L�}����Z�L�h� �[�猞���v�)�BҺ�)�|�$:��Th���0��Y�b��Cpı��!�`�(i3!�`�(i3��Y�H~ XL@3~�����Q_K�W�A���n_�������)��t��?�hV���.�����_ZPV��L�%!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{q��#�i+����Ó�%���d��Gȵ��$6�8(<�����8��	͂'�)�����L��Վa!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��~��ɳ�GV��)�m��G-�#V�"����vg��i<�?���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3rz��G�;����A=&�������9��7�_��ʋ�И_�֠�+��7e���ss�#�-�p��>Uv���ߓD+���4Y!�`�(i3!�`�(i3!�`�(i3�g/t��5�Y�n!�ƪU�\HU���5ߧE4��Fi��|�3;c�<���B�����h�:OJ�R?�6��'�|,kW�A��ˮ��V�rsSRą,LT��ي'�b����|/���d}��[�ƭM�AF�J��f�;�>)�2]MRH�,���
�yJBjbkAޚN��˔Qz��)�3�R�>~qO�P��d��W4���܂�U�ӿt�_ ��N%�Z�U��c-a(􆿳��o ���L�'��*�!N�'�y�G