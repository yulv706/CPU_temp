��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-@���rahZ����*��:�>2/}nQ.��;�p� .��I��u�����c^�.���&��U�,<6V�/���i��?GQ�.��V��?oj�q��8}��	D���o ��Z�� �s�1c��K��ĘV�Z�~����p�l��?��R����lf-[W���f$�J�5��D:mb�@XNQT3�,�?F��3|�N4�����S �n/rq!�t�=�ohWt�_a�7|^���
��0���sW���IᡃEe!�`�(i38�I+�{�Ӓ���h����(Y��h_07��V��&|6�łZ��0y<j]��H]xGMG�2�3�0UhN%ׄ�ns6������y�2)��(p2p)'�8ϳ	}�e!��������߰��͠>��_���t��jo�eW-��ӓ'�al��paf��pD��<��3Z�a�²���C�V�^�"��J�"�퀢W�����*ú��ƞ�qx���J���֤X�j,Zs������gFUB;yB���x	�&"=G�H�D��Lh�&��?N�����Q���qa�EuK�}w�*�*���d����C1zh���
�]S:ֻ�K6ή-��8�#ohWt�_a�k�Ԧhg���'�al��p���B]5)�'�r��'q3�]qLC"{p�G��<��i�m���5�<��~A㉙��[6�)�}��K��;�/O�5'KL[���/*z+d�B�f��!�_��Ҿ��?�4�ʗ�m���;�L|�1��?�1˃�J\wu��v�<f)��,�c�|k�J��-�Y=�#��^ ���L�Y&ׇӭ��h��в���'͍�h\y ˊ�YN��{no�U��^*hrY���F1xH�#�rU҃��~��cC��O�-��8�� �k�IkY�G�
��L�矤�t:(�uO�v���S[W���;\=�H��CW\o6LԪ�u#7z�� Iô͚X?�o>�j��^ :��$q��mKx"E&��� ��l$�������-VLV,Z���ް��!����ˍ!`�^uf8�i�VK9�{F&�z��Iښ��}�2OŘ�C}���\�4�ʈK ������=�����Y�ۻp��@4�+h�	��ދ�*w��H�D�cBP���N�8�c�J���a\Y�����e��rט�������@Ő��t2(;����q�����d�0�YĊ���[ �����
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.��v'gn���1�/�Δ��IgPgud�����`UNP�V��o5]�t���Zu�Ì�s��X�e��ښ�s���I���b�⪒��S �=�[T�)�����5�VY(������b�Kzb�d&(C�#�7#^�Vn���4]�sV�"$�dg�ݚ�Н�:��9KmjWOPg��&yy�;�i*�f`�o�${U��w�X�|0����?�-� 
�FܔR'�Ϟ�Fa��ƙ�Q;��IjWOPg��&yy���͵���ݧG �ŴP��Cn�CIEn4];ˍH���]&�H�ݚ�Н�j}��ރ�	p���{S�GcS�)37J*u��l�M�� �3�~� ��!n}y���q���U��	�,�u��|��].��'���Xw�Bx;�8����*���]�!��0M�p�k�C���� ���:�W@�]�!����=o'Oؒ�b܉����2�V`� �ҋX����@�ڗe'?�<O������9�dMbZ鎬�������(����T�3,�t_-Z��T�\ ���0�:�&^�_Q������jr���~�Z鎬�����;L�=Q/����p��	�ا�*A��]�!��	Ǹ�y85�Q��%s�@�zl���yp��HM�e��`y���MP:��k�_���&:�l�5����-�5�H�^�l��z$
|t�ҋX����{��}��^�w(�M9�5���$����q�h���h����"t��D�e�ȼJzr����x�!����	���q�����h=�%�v�x��*���MC�Z鎬����(S��\� Q���y��Td�#T" �RA9�A
�:��p��mX5�CN�=�s�@"-� �߳G!��1ta7�TD���rs�i�kۜ��/�XO��['���������Y,0=]^	�&������AKd��y c�yO�6i��(�
t��Y�{'%s=ͱu��̦�"�K�b��Ub�ۙD^�V]��}R�wX���o�K���d7Ud䙌�!�!7��TD���rs�i�V�W�+1M�`�"�X��O�'{�,0=]^	�&������<y�׀%\ʞ�sB�_�6�vg;Je'���Xw�!�Tcִ��#"�餯���Z鎬����l��f>��d�����N���qH�iQ��e�Z鎬�����;L�=Q!s"֛
.C���~���J����m��w���Z鎬�������(����T�3,�t_-Z��T�\ ����`���Gé�ĻP�q����0��9��?I��w��,c�A�L'�H�N�P]��Z���Ga(􆿳�b�툛�*�}r�HDʞ�sB�_�	�/��TD���9�,�w}J�A�D�Q,��,��u����	a���*Ѐ��&~�>P�2-i_���F��.g��4������	a����DY���%�a��E=��}�У7ְU��d�٣��c�A�L')6�Y������i�t_-Z��T�\ ��9O���t�6|z�ä�@�i�f�UY�h�k/���Z���{lIk`��L��s7s�9���o��S8�'�X4�B�F\���e�Qi��S쑧��8���/�l|�*"k��c��*��#�|.�Tӏ+~'%�ͫ ���X��֑xGV�z؝s7s�9���o��S8��I
�R�W4�b��nw;��ߪ��w������d�x� �qsC�CW�[��k�6o��d�٣�����6>���3e���;�/���jbPh�e�z��;��]�!���1����mZ�M�R���'�r��'q#�� �[N0V1�M}��E�]�!���1����m]^U�*�!�3oz�2Y�{'%sgeߪ�{o�${U��w�X�|0��9)�����m��/�	1I�5�e`��9�'�E�Jg�LA�dWH�:�g�"I7s�9���oC�M��N�۶E ����C���� �u|Z�x��f�=���Z鎬������Ȥ�8��V,Z����jC ��+�Og����n�e47�O�T��ڏ�j�j]��n�hy@k�.�r��V����*hq5�*�,��-��W�v	�KT��;X�'�(+,:��~�Db*��E�&����f��jvr��Q������h����@$˺/t��꫕qŧo��K�O���J�Z�@^��}�/����p��ey�u���FR6ni�N Aj�]Y�{���O&�s�N?5�ֵC8'mX���nOU)���� �Q�c�C;=B>��ʅ�<��W5���!Vi��%�e�TUݧG �ŴP��CnxPT����L��S7-�;��|B* ^���x��A$�P�De��5�B�7Ū�v�>mW[�Ƶ\�����Y;�I��c-(��nr`+� ����)c N��r*�Ã�mH9��0�zG��x{^4��*mxMV5��6_j��r�.u|Z�x��g����ҍ�f;[���=�	�:˳����
�?<��{
��>��Ǉ�y��s��U;4D�f�b�Hwz��c� �@w���H��j�Ï��	�M��.�X�3�� �f���=����8,b���-M�O��~�xMV5��6_j��r�.u|Z�x��g����ҍ�9g�M�G�n f�Lu�m���������f�iC������t�f����pD��^A��xB <��g�^&����1�A�O����L�7��3�/gWaU �Ia�<d��d�J/�#{�mW[�Ƶ\� �Ģ��|�-M�O��~�?Ohk���0La������t�f����pD��=�<�^p�-a�D͢q��`�L. � s��/���jbPh �Ģ��|�-M�O��~Ӵ/V�S���/���jbPhŋ~���%.�$!q��)�'٥��gV�J�1��씑�:��KY׏�����Mrw�&�z<aSm�6��`4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY����|u��IX0F�M��܉=�!U��s��'Y����]�Y
L�1�'�E�Jg�R����+�AMm?��%o�w���iqI�����I�d�`��L��s��It�Dʷ'�r��'qm�±��m|H>=tL_�+�AMm?��(xʶ���զ�[#�Qf�'�r��'q#�� �[N0��r5v��|�
9g�M�G�n f�Lu�mz���5|���;��Ѧ��c-(��ܬ��x��!_���{� ��b�FP&���g�|R��q�g���c&,�U������v�sk�Tm�k]m��7s�9���o��S8��Kq2�譾b��nw;��ߪ��w��f-�&B�����v�Xc��m�)YC-�T^*7s�9���o��S8�5|���r�\���e�Q�mƿ�Lg�g��U-�e��C- ��b�FP&�I�_Pg<����v%��cZ鎬�������(���-y�5Y8' �*�I��p��HM�e�Nu�5=��{=J������P:����\�W�EC�2[QvA�#���?�Z鎬�������(����CCю�l0�7��65��Wǖg3�MM
��,=���L�E����L������Jn,���`&,�U������v�S�w�KIOִ��#"���L��ǿZ鎬�����A�p'�:���=Aϔ�<"(ZW��ό���.ӌ+U�HJ�h<����y �h�6Q�7�ǃ4j�mrY�{'%s2�ew��e�X�+� �{�c�vI�ߪ��w������g#��� t+mm� �8���-�r�MM�6�y#�c$?��ό���.ӌ+U�HJ�h�����|��Km�^6*�d7Ud��_Y1��X�#�c$?��ό���.�B� ��~���1`|5��[&�$*�9U�&�(���D��N�j�W���LM���9�j)�����R���M^.��	�+|VO�⅘�dN�<@Iv���a_|�����	�͆�C�_]FP?$�N(p����c3ჭ?�\���3cx���K*F��}v�R"l|�*"k��͆�Wu"���S���Msc	�ۮ�|M�U��(p����c3�C6�=�����!���&v4�<0�����R�Ӥ�D9w�tkb��u�"�^���9f�vr2�����C�6��{<v�/���jbPhM�x���I�c�Z�~ɞJ$��^�5M�YYroE�4rh��|��3���ʪf;[����h�����#8Ԧ�/�w`�e��>|z�ä�@�Z��&61��7LF��4�֧��L�q���Ᵽ��E��dN�<@Iv���a_|���?��Y}��d�����N���qHTZ_&bq�f;[���0=�!�hj���*6S�4��?��kR�KC�m��Of�!���ٸ���<�ྫྷ��c\?
������'DV���8Fv7˨�c3ჯ4D���t���\@'�^����t���3�l�^s�kQ��b~*��s�F�KD�Vr[/}>5��0*�ߑ���7��3�/g�d��8���bp�a��N}9�˕��76�>WԆ.l�I���{�IX��WG ��d]��>���}r�HDʞ�sB�_ە|����<5��H�3-nmW[�Ƶ\�ŋ~���%.��8;b��U�����W���c-(��ܬ��x��!�GE�i��P����{�/���jbPhi�x�X�a
"xT��z�����~ԑ{�χI@���̎��#p��T���ڙ(mY�����È�Fe9�\�W�EC�2[QvA��>�q��J��ΥT�t-}ʙLY�>U%����f�4D����G9�:Q���i�֒�B���5n�[�f���r���˃�I�H�Nb�*Z鎬�������(���o�HT蔊��8C�\�`��L��s-�aS6�0�7��65�����S3N8BW�R7���r_��mg֓:lla�v�r���f;[��སf�B��IȘ�i�E�����
�?<�v1a{J��`��Ks���ɛ�?ө�h�����#8Ԧ�/j���྽P�\�2���?-Sah�/�����ྫྷ��c\?
�����$�,��wZ���{lIk`��L��s���:��KY׏�����M�}�u�0�_!�`�(i3�K:+>5��H�3-nmW[�Ƶ\�ŋ~���%.��8;b��U�����W���c-(��ܬ��x��!�GE�i��P����{�/���jbPhi�x�X�a
a%��w�VW���cl�����<�������=�<�^�
E�4.��̓u�J� f�Lu�m�k]m��4D����'٥��gV�a�;�f��h�6Q�7������w�j�W���?E�!$6������1g�W8]��?�̟�1�+�9-�i"'���Xw�j�7�� [��ѮT�<��{Y�7k\��ϡ	t$���!���zl���y(ɹ�f=�>je`��@d:�����{~\�e�E���Q'�z�Mv!���xL�2�r��Km�^6*�d7Ud��_Y1��X�Jh�o�p��Hp9��Ǧ"�7�F�Q�Y ��b�� 4��P�!�c�dN��B���t^deZ���{lIk`��L��s�Y*&m1/��f���r8,}'�%�y�P�HS|�4�04�jfJ�1����9�8;}P�%bGq��7ʶ^��v$���D�<D��-��r��}m�]9qI/��\]�S���M��G#��Ll(��?��kR�KC�m��O���nk�b*�����1"N.5$R��
�[b%Ɨ�G#��Ll(��?��kR�KC�m��Ob�� 4���\�W�EC�2[QvA���]F^�	rw�&�z<al����HZ�D�$0�	W��^$k�6P�p�HZq�A��Д�TKݚ����0��s��@^��}�/����p��M��R^�h�0aQ���A%z�X�*63�o��a03��(�0��x��y�o�P�~�����*�����1"�(���(p����c3��O(����8+f«L�I�_Pg<�ZVv ?J����xK�h�6Q�7��ҿ�Gz���D��B�UX���e��}r�HDʞ�sB�_�����C�&����1��Νg��$/���jbPh���ʼ�D�u�t���Y���I�9@'n>�I��Z���{lIk`��L��s�x��y�o�P�~�����*�����1"�(���(p����c3��O(����8+f«L�I�_Pg<˙Y�#�{U�xMV5��6ִ��#"�BcRf`�B��ΥT�tɞJ$��^�5M�YYroEΖ�1�!�fC6�=�����!���ԓ;(���[b%Ɨ��O(����8+f«L�I�_Pg<˙Y�#�{U��D����'YC-�T^*������YC-�T^*�����5Ou�>����9��0Y d��4D�����p����8z�mx�ݫu��w��a�%�Hw�<��'&g��h��P�l��vE7�MW�}r�HDʞ�sB�_�����U�8BW�R7���r_��m�%&^�nƒg�|R��q�bĬ؈��0Q���g�����bo�P�HS|�4�04�jfJ�1����9�8;Hu[[Zq�,�%�Yo:#WQU%����f����gsN�ސ���*���mЎa�<d��M���yt7�n>�I��Z���{lIk`��L��s�5l��['P�!�c�y�&S��n�Ut�\��Msc	�ۮ�|M�U��(p����c3�T۳�͕���D�$0�	W��^$k�6P�p�HZq�A��Д�TKݚ��91+�Z��5l��['P�!�c���px��=n
V~$��t��i�4W'�*7J`S��H��efm�0z�cULPz��E���"�K�b��Ub�ۙD�X�:�{��>je`��@d:�����{~/֐��̺���<���#�x4v�mw�xȀ��D׏�����Mp�-a�D͢q��`�L��˓#����Msc	�ۮ�|M�U��(p����c3��5ߧE4��Ћ�E?�B�n���5�����
�?<��{
��>N�q"b��C��R�f%�.(�q�,k!��L}Y<� �ѽ.�'�[�b~*��s����g�|R��qj�֎���4b�-fz^�	�ZXĒ*C���� ���ۀa���n��뾦����pP�*���k�<_^���C�Zҝ;�+�pʷ���Ϡ��,�%�Y�BI�yא]`�"�X��O�'{��9�]Z-�[�^�o�R�1m�I�
Z�9�d�L��!�&�4_]F�Z��g�d��%�z�J��=�	�:˳����
�?<s��WM����x�ԉ�>�"L?��� e8�~��	W��^$k�6P�p�HZ~�똕<�/���jbPh79 ��/6�tTi���׏�����M>je`��@d:�����{~�4�%���J����Y04t�C�"���z8+?� e8�~��o:#WQU%����f�<���Hn
V~$~��є27�C���� ���ۀa���n��뾦� e8�~����˓#���~��є27�C���� ���ۀa���u�1��s f�Lu�m�c5��3t���=�4�04�jf>je`��@d:�����{~=�	�:˳����
�?<���z`��k��f�iC���B�_�+�)#P�j2E�?x(�i��/R�xȀ��D׏�����M���pP�9��0'����f�iC���B�_�+�)��h;�ab���c-(���dI�� �p�-a�D͢q��`�L�5ߧE4�� �U�O��. � s��/���jbPhi�x�X�a
0��d�����ސ�����H�^W3����4��ܧ4��D8�>=�o*�F�Z���1ǺvK}��a-6�Da�\�"7�D�'٥��gV�T۳�͕�𐮋�Y  ��!���#k�˟ܒ�o|k�Lb�~������VR��)Đ��hJ�L��Z��kM�8�"�^���9f�vr2�d��-��!h�}�M�����VPYUt�\��%&^�nƒg�|R��qưb�����|	ҷKD��x�ԉ�>��˓#���0���7�0>�Q�k^�ïw��O�$FP��{�/aC6�=�����!���P��
���j5�/?:��5ߧE4�� ���M�����.b���-��qs�VY��bE�^2`�"�X��Nݲ���+X��WG ��{�χI@�괆���-VL�[8�[Kh8,}'�%�y&����1�^M��C�\	��rR�oʒ�^����V�R+����KVY��a-6�Da��yU\��À_)WG9�:Q���i�֒�B�B�R���>_���d2<��k]m���Wa�>�q��k]m��z�q�T�Ƴ8,}'�%�y#k�˟ܒ�o|k�Lb�~������B�fL�ŏ��Sߓ�\�)�w
��-M�O��~�-}ʙLY�>0Q���g���C1zh9�n�p8�#,����C�_]�#}h�[b%Ɨ���7LF��4�֧��L�q���Ᵽ��E��w����F�'�r��'qm�±��m|4��+$#k�˟ܒ�o|k�Lb�~�������oF�t!�0xޚm[Ut�\�����駈&����<���՞e{f�!���ٸ��.�[ ٓ��r_��m^�=�L�v_����xQ�n
V~$`;��@�+;�6����O���H��`��Ks���x�ԉ�>T۳�͕���CnX�&��v~�z�xE�?F ����4D�����Mv!���xJ�1���)�@����p�-a�D͢q��`�Lt���3�l�^s�kQ��b~*��s�F�KD�Vr[/}>5��0*�ߑ���7��3�/gWaU �I��z��R�C��%�!�uV�Q���a-6�Da���1j|g[Ҡ(Y�u�o���z!�l�P��,J��La������t�f��U�~�{k���!q�����
�?<��{
��>�&9�`��ͧ�˓#����Iw���L�8���-�r�MM�6�yJh�o�p�+���8�׏�����MJ�1���ظ����05 S�s�l��yU\���i�֒�B���|��j_H��;Cj��a-�a� L�/�{.;2I���;�XNt~e�1���'.5B�L'��:�<X��u�>j�V����%�>.}2�X>�Q�k^��vZ� �/Q(�?�\���3cx���K*F05 S�s�l�?�\���3cx���K*F��}v�R"g�y�ޥ-j����*��Z�ࢸN��_��+��d�C����13�3��ŧ���X� 7���s'F�j�W���?E�!$6ӷ:���N3!GjW\nVU�NtZ��\���Jw��3�ɞJ$��^�5M�YYroE�4rh��|���'��<���XQ �Kk�2�:,crۈ�L�o�!�0Q���g���C1zhi�Y
�,�ӎ�Xp�,4�֧��L�q����*Y�Pܞ\^�5~Dy_���W�>y�۠����(kp�~ge?���W�>y�۠����(k�pS�yW� ��푮1�r^M��C�\	��rR�c�3'A��0�7��65���KVY4n8�%�(%�ɏ�X,���֑xGV�05 S�s�l�?�\���3cx���K*F��}v�R"��s��U;4^M��C�\	��rR�oʒ�^����V�R+����KVY4n8�%�(%�ɏ�X,���֑xGV�05 S�s�lrn�U_����m����s��U;4Vq͜G�Ɂ�I*�?��m�±��m|������E��� �r#�j�����'J�����d7Ud��_Y1��X������K׏�����M=0�&ǧ�"�0K߸��S�Ȍ�>>Y�k9;��|B`���m�Q�@��߿�܂��I���J��<��%�8�cqQ��ح(���|�ط�64[`������r���aM"���Ig�{	#YHN�����Z���삕��y��}�p���P~����F�9g�M�G�n f�Lu�m��jЏ�_� f�Lu�mQ����`��'C�>��/����p��BZ��L(�0Q���g���C1zh9�n�p8hѶ���� f�Lu�m�� ���~�0Q���g
3K�������: a�`7�H'` �#�W����;���EWrC6�=�����!���w��z䮃������4oQW*�dsk�Tm�k]m��7s�9���o��S8��Kq2�譾b��nw;��ߪ��w��f-�&B��ZӔ	�2��a8´�*�����1"�H>+�w��0z�cULhv�R�+Z`�"�X���!y(~,�a(􆿳���/�	1I��+U�HJ�h60�,C�����-VL�d�٣��c�A�L'�ћ~�i����Q;��I�t_-Z��T�\ ������W�^(�;���EWr�?�\���3cx���K*F��}v�R"7s�9���o��S8�i�۲da�`�"�X���!y(~,�a(􆿳���k�H�H�g#���MΡ�@�������]�!��v$�7<� ��b�FP&9g�M�G�n������#�c$?��ό���.��4oQW*�dy���jl7s�9���o@�ڗe'�g#����t|Ơ$��#8Ԧ�/#�c$?���rs�i���%��v���0�BE�9Y}��P���"X��[�`�L�iֱg#��� t+mm� �8���-�r�MM�6�y#�c$?��ό���.��4oQW*�d�Y��>%��Ș�i�E�����
�?<�v1a{J�ǃ4j�mr�q���U��.hU�����x<��z���76k����9E-M�O��~���
-m/�k]m��l|�*"k��͆�Wu"�z�X
3kZ��z�������omi7x��8fDd=ܙ`	���d2<��k]m��l|�*"k��͆�Wu"�z�X
3kZ�?�\���3cx���K*F��}v�R"l|�*"k��͆�Wu"���s���刜t��i�4~f�@�f���j)�����R���ɞJ$��^�5M�YYroEΖ�1�!�f�Mv!���xőT�ZS���c�Z�~xMV5��6ִ��#"�BcRf`�Bf;[�������v�� f�Lu�m̝' gi���Mv!���x0���7�0>�Q�k^�ïw��O�$FP��{�/a�Mv!���x�h�����#8Ԧ�/�w`�e��>|z�ä�@�Z��&61�>����'�r��'qm�±��m|/�l�`�Ђ�nF���]�Hlu���"����r�[O��ɔ�<5���3��< ���m�QA�Q* �
E�4.��̓u�J� f�Lu�m�k]m��4D�����Mv!���x�}?�N�*����4����Bf����{_8�Y�����ƿL?(��^9[�_Q�������3���ʪ��ΥT�t�\�G���(?"��W����_�M86\�4�@����s��X��WG ���05/������3 ����76�>WԆ.l�I���{�IX��WG ���D�$0�C6�=�����!���N�q"b��C	��Z��5�_j��r�.�`�u�?ϗ6�+b�f� f�Lu�mj��1�-��h9x�����
�?<�N�jH'�7<(�lb�<�䛄��g֓:lla�v�r��ɲ�ΥT�t�
E�4.��̓u�J� f�Lu�m�k]m��4D����'٥��gV�-}ʙLY�>U%����f�4D����G9�:Q���i�֒�B���t^deZ���{lIk`��L��s��9�W�"7�cL���	Ǹ�y85����NZ �~�P��?
������o�ؕ a�o�${U��w�X�|0��r1U�%G����pP�h�Qf�\�e�E���Q'�z�Mv!���x��f�B��IȘ�i�E�����
�?<�v1a{J��`��Ks���ɛ�?өa�;�f��h�6Q�7���O\f������ �r#d��@#�h�Qf��	y��J���gtb4�^�q_ϑ{�ș�@^��}�/����p��\�<���+J�1��씑�:��KY8aw���`f�k�X��0�/�M۴� ��h�6Q�7�W-)Վ7�t!����}_��f�iC���(b�Y6F9j�7�����C���� �D,��a��gWaU �I����~ԑ���d2<�U%����f������U�h�Qf�fY�J�]�d(����D��Z�خ-�D��~4p��T�����Xaw,��� �r#�j�����'����v�?MN*����h�Qf��	y��J���gtb4�^��r\�����H��efm�0z�cUL���6磌^�|U߳��َ��7�np���� ժ��[:0�7��65�����S3N�xȀ��D�[b%Ɨ�{�χI@���̎��#m�QA�Q* ���h�����7ʶ^��v$���D�<D��-��r� DS�
��c�Z�~��$�����P�\�2����`jS-Y1�b�o��#8Ԧ�/O-�4'h������1g�W8]��?�̟�1��H�^W3����4��� {�'#��c�}���Fo|k�LbJ�1���)�@�����9�d�L��%�2X��<�(xʶ���aG���z䮆G�_02�����W\D��	y��J���gtb4�^��EB�?��ސ�����@�`�\�e�E�~*�<�[�4b�-fz^�3��(��w��a�%L�`���žj)�����R�����
-m/�k]m���Wa�>�q��k]m�������5OxMV5��6ִ��#"�BcRf`�B��ΥT�td�4�t��Է'�r��'q��{����f;[�����a�z6�>��M\p�� f�Lu�m�=n$��,��5�Q� ��5�gZ�W���s3g�W8]��?1r����X��WG ���D����'YC-�T^*l|�*"k��͆�Wu"�z�X
3kZ��O(����8+f«L�I�_Pg<˙Y�#�{U�?Ohk���0����*��&�Hx��_�=�<�^�����x�����Xf ��zR��%�>.}2�X>�Q�k^��vZ� �/Q(B�R���>_�@���J����p���$�J����3QP�B�=s������m%�td7��|�����ob.�Y�2W����xK<y�׀%\������Jh�o�p�Dՠ F!5���٠F�]؇��k�ঢ়�?{���X+:�J�oСJb�C$�-���}r�HDʞ�sB�_�����U��xȀ��D�[b%Ɨ�ɞJ$��^�5M�YYroEΖ�1�!�fC6�=�����!����&�q?Yx(�i��/R�P�HS|�4�04�jf�,�%�Y�iw�|�ݭ�̓u�J� f�Lu�m�k]m��?�qjv
Kð��T�ҍ緫ĭ?�\���3cx���K*F��}v�R"������YC-�T^*���:��KY�[b%Ɨ��o�K���d7Ud��_Y1��X�j����v$���D�<D��-��r{R�@Mvc�}���Fo|k�Lb_N���9���VW���cl*���k�<��~"3B�>�����3����@ 0aQ����p*��vE7�MWM���yt7�n>�I��Z���{lIk`��L��s�5l��['P�!�c�y�&S��n�Ut�\��9��xe˰M{�?I|z�ä�@�Z��&61�"L?��ٶC$�-���0o��,� f�Lu�m�=n$�4�	t�ܐ�ސ�����@�`�\�e�E�~*�<�[��x��y�o� e8�~���ސ����H�Nb�*Z鎬�������(���fx ԣ��0�7��65�ⲺŜ2mz�X
3kZ�B�R���>_M��ZLh-�� ���$�� ��6A��e-x�_�3t���=�4�04�jfp�-a�D͢q��`�LT۳�͕����t��i�4~f�@�f���j)�����R���rw�&�z<a�i���i��|:w��!C���� ��`�u�?ϗF3t
��
������F ��c�ϩ8{8��d}���d�d��-��!�j���]5M�YYroE:�k*�.�mo%��`���a-6�Da6UQ�㔩�(xʶ����y5}�E�Ǥ�Hp9�����F��;�D�$0���Q8� Lڈ�|�<���H-�ȎBu�h�Qf��!yX[�C����i������^`�|��K�z��KVY�/̥@X�4�D�$0�\�e�E�0Hl&p?�ð��Th�Qf�=�	�:˳����
�?<s��WM����x�ԉ�>���pP�h�Qf�=�	�:˳����
�?<���z`��k��f�iC���B�_�+�)#P�j2E�?J�1���#P�j2E�?T۳�͕����L�ΪA��VR��)Đb'�Y@%�F~ʽ�Wn
V~$��L�ΪA�ʴ�!ޭđļw-b�&�I/��\]��a-6�Da�/V�S���/���jbPhM�x���I�=�<�^ e8�~����˓#�����9V�S^��f�iC���B�_�+�)��h;�ab���c-(���dI�� � e8�~���5ߧE4�� e8�~����˓#���~��є27�C���� ���ۀa���u�1��s f�Lu�m�c5��3t���=�4�04�jfc�}���Fo|k�Lb�"L?�����9V�S^��f�iC���B�_�+�)��h;�ab���c-(���dI�� �c�}���Fo|k�LbJ�1���)�@�����9�d�L��%�2X��<�(xʶ���,������P�>|w!&&_[j�/ྫྷ��c\?
�����_U��A�3P�!�c��j$���-M�O��~�Y&jV��hK��aF?����:��KY�[b%Ɨ�őT�ZS��A��H��c�}���Fo|k�Lb�05/�����VذQ��k]m��
�HYF�@�9g�M�G�n������[Tj�qM�3�HK�zV�v'#`�x��X��WG ��d�4�t��Է'�r��'q#�� �[N0G��0n��ƿ=�<�^���pP�vE7�MW�}r�HDʞ�sB�_��F�İ��|���T��(���XQ �Kk�2�:,crۉP�HS|��� +\�?�����V������.b���-��qs�VY��bE�^2`�"�X��Nݲ���+X��WG �����d2<��k]m��������YC-�T^*���:��KYD@��� V�g���ޔ[�,n�v��"q���^�o�R�n
V~${�χI@�괆���-VL����v�?MN*����8BW�R7���r_��m��"�oi�8+f«L�I�_Pg<�!�V�UCb�z����8�@ؾ�X�rw�&�z<a��r����K:+>�B�fL�ŏ��Sߓ�\�)�w
��-M�O��~�,�\����J���o3c�-��;���֤���n���v���=�W�� ����:+FwaT۳�͕��-}ʙLY�>0Q���g���C1zh9�n�p8���$y�J���o3c�-��;���֤���n�j5�/?:�x(�i��/R�-%��ʦ0�D�$0�ސ���9��\��E��%�z�J�����1j|g[Ҡ(Y�u�o���z!�l�����C�8BW�R7���r_��m5%�h����v'#`�x��X��WG ���S�V�C�d�����N���qHTZ_&bq���ΥT�t���pP�h�Qf����1j|g[Ҡ(Y�u�o���z!�l�����C��xȀ��D׏�����M����V���rw�&�z<a��r����-%��ʦ0rw�&�z<aIP&_V�t>�3�eZ~h�����p�S�CП�_��r<+��Z۳
0.{�R�$�V�J\X����9H\WC,���Sߓ�\��������\�:@�8�xMV5��6�Y^8������.�'��}r�HDʞ�sB�_E�Xf}}��v$���D�<D��-��rv�V����v$���D�<D��-��r{R�@MvxMV5��6ִ��#"�h�6sՑ����*��4����QM@��e]����X� 7���s'F�j�W���?E�!$6�AKd��y c�󐪽�r���8��9�8,}'�%�y�	�ؽ�3���XQ �Kk�2��Z��%v���}r�HDʞ�sB�_��F�İ��8�7��0��
! R�7��1�G�Qc�k]m����\[���0Q���g���C1zh9�n�p8��U��N�`;��@�+;�6����Y�-�_{sx��)�p��6����O���H�Ԧ)�,�|^�Ő��ngL��k��TA�l�Lɼ�wj���P��zl���yf�^S�l��*s���j%�ɏ�X,���֑xGV�05 S�s�l�?�\���3cx���K*F��}v�R"��.�[ ٓ��4]a�#�b��nw;��-�?I�g��Q;��I�@�����Ut�\�cI��S}H-��;��>�3�eZ~-Y1�b�o��#8Ԧ�/O-�4'h���˓#���0/zﴚ�:�L�������-VL\�806����h�6Q�7�8��x$�v$���D�<D��-��r{R�@Mvp�-a�D͢����3�$Ηw��S35�����߸��S�Ȍ���#�X�6j�"Hs[Y��N(?a5���!Vik4�݄e�k��m6[��e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@�ޗ9(����	�^��i�{���_�-h|,���(����>S��ә�����/�4�}n'���a*�x���� ��V�h����� ��?)��h�dZ�c��ǌM̯� VU+I���ť1k�`d��q�G����p��=.,����k����씧;�y������,�p���>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z��r9�3/�OP�I^���V� D;5B5Y+�T�����N�܋�z2��~����ܷ|�p�6 �P�{n�da*;��;ۂ��IÙ=�H(c]9禩�5�Y�w��n	~����=��q�a\Y����_�G��GJHn��z���Z�n����t���i�Oa�b׉�^9Y�rU��6���h��J�1,!��a\Y����_�G��GJHn��z���YG�sT�Ș�TDв�0Z�׉�^9Y�rU��6���h�X��-�`V-u9�`�JHn��z���YG�s����Ӭ�oi�Oa�b�����I����ʮ�&3�-��_'��-d�Ry��\�v�[������ڶ�!!�+�R�G�Qr	�%\*��t���Y
 ����6?L���^ֻ����XP����d�ӓ
(~F�iO	������9`�p�0�B~W�u���iL�&Ш%� MjCЭ�J�1,!���i=���[&��?��
JHn��z���YG�s��K������-w˕��F��v_}*�����i��!�����9���k��h�@�sj|~��A�!`�u�!j;5B5Y+��q	k���Ak�$����v7�'��O�q�Yz��"�ձ[%�U��Q�f�!�+��7P��T�<��z��}�צ:�)��-��7�Sc�Q��~�z��e�K����{l�f|����%Hlܾ�zx�8���#�!� k&oA�\ֆ-�֥�� ���Ig`i�ҋX����0�a1i~J�5�#(�@�%PX��n&oA�\ֆa��M(��E��jh�m!��ʧ�9�x�^4/��?Ev�~������]�!���R�qSe4�uS�4q�
��n��7��!n}y���q���U�M\R�'�k�!!ʽ��n��7��!n}y���q���U��֎)A=�s��]b_3#ڸZ鎬����8�������F�!���Fi����o_3#ڸZ鎬�������l�T�|�1��?���HEcx������]�!��	Ǹ�y85�:V�Fx��Wǖg3ȓ8���/��x�����^�o�AZ�Xh�c�Q�j+�B��oy�{��vvfۛ�
�B������;�
�{�L�t��n�|��].��'���Xwd�n]N����=;���Wǖg3ȓ8���/��������,J�l�/�E�,�h#Q�?��}�1+��%w�[�O�r�CC��5��y0և��@�)#��O��t{��*�cw�5>��Г����1���I*�?��m�±��m|i��%H�	S�)37J*uc�A�L'�t�N)�~T-��qs�VY���/7R�%�T�\ ��a4�0 o)�J���o3c�-��;�����!�!7�<��z��}�0z�cUL�JJ�4(o�a\Y�����BT�^��a(􆿳�b�툛�*�}r�HDʞ�sB�_�	�/�<��z��}拋ġC��ױ����h=a����gW��_K����(�
t��Y�{'%s�O��W��[�$��X�l�Lɼ�,0=]^	�&�����虭Og?6�������O��X��M�TD���rs�i�ק)"�僁Զ$�H� �b��nw;�X��������`y���M\R�'��5D��0h\Ef�>yf��i��]�!��$��lW�d&�(2���7>	�����T�3��]v��#�(ic Oag�qod�֓�����p��=.,����k����씧��a,�>+�'�.�P�I<���V�iC�<�Vz���@9��P����eR����i� �߰a�P�Fpwi�����\�v�&��sf��`�|��K�z������u��C��J�hx��W�D�U�6g!�Mn�g�?Q��G���@Ő��t�xU:풲�>�������K�QB�f�%�+I��=Y��_��ġC���&O�ǻ����������Cos��ǉ8�!��Z��beNY�����$#Z�����t2FSx�lޞ�ό���.���K�Q�t���(�x��V��ⱹ�(O,[ǘq���U�pzl��a��&5�/h�t���(�x�/����d�٣�����6>��b02�O �+s�ɔ��]����ڙ1�ٽ�H	�]�!��s���X*���Zr�lR�����i�}��Y!��]�!���1����m�6/z��:�	Ra�v��E+����Z鎬����Y�V��#qˢ���[@;��o`��G��]_$��=Y��_��ġC�����K�Q��L�
���=�\[L�ﻋ-�����S8�F�Z!���{:������q��WX��y�g��U-�e5��e6²�n�\l����mAp[B�����'���Xwa'�<� \:h�����ի�~����q�
�Z鎬����Z��C�Ջ���`���<��r)3<Wu|����d�٣��c�A�L'D�j�b�A$`�y��������\jt
�ߴm�R�wX����K�Q��&���S=f�?TY�͈9�4�Րﻋ-�����S8�qT�8>��ڧZ��7����.C̠�&A���T�\ ���|.�Tӏ�٪DX��1�gB�� o� c �_�K��ՃZ鎬����Y�V��#qˢ���[�'��O�c��M]l]�F7�Ghjg9��G�.'���Xwa'�<� \T
�ߜ-��ِmd���u�a��b�hΤ�`�ό���.���K�Q����/�4O�#��K��%r]�Bа"�����d�٣�����6>���ZLl�]�̑�z����.j�l�&�ﻋ-���C�M��N��+w�7�.�@��>�̑�z����.j�l�&�ﻋ-���C�M��N���<n��nN,�P-��2�|�I�7Sx�lޞ�ό���.���K�Q�P��G�"�]/�����:�^��ר:9f��c'���Xwa'�<� \�]VI��Z�v��#K�ϩ�E�m�ﻋ-���C�M��N��|�F7�_����'��e��"���N�@G�"Q��'���Xwa'�<� \%5�Ψa����g�cЉ�M��'ˑ�sO�rs�i�>�Ca��?�o>�E]�٩��7�v�ԯ�z�C���+w�7���\(FK��WdM4@Ȍ[PP�\��]�!��	Ǹ�y85�ٙ�횔6�a\Y�����BT�^��a(􆿳���Qs�����T~}���`Z����<Z.َ��)(�w�j�d�٣�����6>��b02�O �+s�ɔ�7�9���������D�
�ZM��9�]�!���1����mr,��>T��wy�㱏>1�gB�� ��U��#bx�d�٣��.���ᣓ�)�3�#G����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h���[m���~������a����N���#t����n�~����p�@����9)����K�d���tn�u�$d�I�v`J��U����+=����7�>D�c�lQ@��~�
�KT\�mɍw�B�I:׷�F�20)�_SsJjvCn������Y�
���h$�7�R?�6��%]����	����X����(h�š�b)�pU
0
m�k8�5�>�yKYQs��[�|�F��ˮ�pd�Zз���\��6�R�X�?�I��H���Ku U�zjb01
�;��S��y9Ez��}��H֞��� �z��w�����4L"炡t�8j�t�Y�Ij���0E���FZ���;D8���:��M�S�ᳰ��X�z���t���Xo޲G�����$7x�c >��}f]���]�w9"x�g�Hz���!Z�>��P$��j�f��>0M�<k�lw�i}4���0�H^�wr�y[�qj�15���{v��_G.B���uOܟB8�A��jeN�V�������1d��3+'P2ӡ��,����|#^�Vn�B��מ�\P�O����X�e��rl���1)�*C�8���EBy��J�z�3���X�|h���	a��b�u�/�'���j��7�)a���%}D�����!��g�-��\��OA�=�~�]��d�Y��o�6�֟�Zl��9����WI�;�_�	�t쩖NUD60L�b�J��@��y���Y
���^�.;��L�O<^��`Y�F�����I��#��
Mc��������=��:p��C��8�@��y�.��3��pƼ�+2!n`�pάYc:�IX[��O2 7�,�)�C5�!f�f�2�c���w�LnXZh��\����L�Y&8���p�lŕ��W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+�S�AZL�0hs�A_	�K�o[��mU;լ^<���X�E��~d2����eI���%�ׅ2�����Vc2�����Vc2�����Vc��Y7�<�L\��x�f���4/C³������sn����,�2�����Vc2�����Vc2�����Vc�cRq>h$8'h�5NG=���YC�вԺL�9�<�=CFswd� l�\�n!�X�%w�"����e� ���"�t��k�|v�<���5�i��p"�.�^�h�xs�MC�%`z}���6W��k�L>*Ǽ0�&���v��t"�~o�D.�1o��gE���Y"㖹�� �����@����nn����^�o�A�ސ���zZ
�
(ȳ��(��$�t�r���޸Q;�G*p�[��
@נg����}@o��Ӟ���}T����;e.�����$�q��T�G�'
c�����H[��e��U��1(7�����n�Y������ӈ��Ӵ�K7K	Z�ǚU��x�n���y�1���.R���oKL���:�af��pD��ɬc��WN\bE�􀈺� 3�j U2��EE_������i��sRZ�Z��*^QP�o4f��I�A���Z�@�'�B^��T%Ǿ��;�>�k��?��9)��:�����xO-�Y�il�ٙ�}M�32)���έ��2F����ӳ�Y�
�q�^ƩW?�d���&�J�-|+�*��'��e����9��������U���u�\��~��}�P��{�]���q�GR��r#�-m�]����ڙܤ��[�p^����,�ǰH7"LTftTWT0z��c��h.b�POlb�ui�1j(���WV�#a��mJd��?�7r���g��O�?Q�d�:�u��������Ѩ�f?�R������R]Y��5��X@w���H��j�Ï��	j�ە�((Ut�\�5�UI1�gB�� ]�Q%�%��v�ڕ`�c����������'|F��ΥT�tT۳�͕��8j��y�����_��
�Q�Xn8��2�ֈe-M�O��~��D�$0�����/�0k��DyR*E���&�Ut�\��R��13{�]���q�GR���1��X��WG ��c�Zਧ�%̑�z���o�+~KO	�c�Z�~�{�Z՟|
�V��&|6�łZ��0yI�[	ϱϲ�ΥT�t���pP�h�Qf�m��"���@��b�x�. ��#P�j2E�?��b����(K�Tl�;���f�����q9+t�}�xȀ��D׏�����M���pP���._(��O�#��K��%r]�Bа���/��D��c�Z�~c�Zਧ�%̑�z���o�+~KO	�=�<�^p�-a�D͢q��`�L�5ߧE4��rw�&�z<a��N� φ��<�6�Ps_*�Gq�p���xg����6�Zk��E�? ��hID��>��9�=���@	Q����c^�0?�d���&��I&�^��"zQM��7��J��mE0�gǞ��D�r�c��orǟD�ui9�f?Y�O�`�MϦ��pCeu��|̧������$Y�G_Q#j<��#�Z�/�k<����o��Ժ��e�����Ԓ���g���	~���;A���W�>����V;5h���X �Z�^6B����B��E��G���ِmd��
/��y;���W����Dh��Th���X �shf(�`�X�G[��P�'�h�&g?	��o���E)��k���I�w�Q?�y�"�]����ڙ�k����ˇ���������76S=f�?TY�ސ�����)G�J�cbp��'@
9��y��%��3��ןmnRYpW����@	Qq��=��$Y�G_Q#j<��#���z4�����i=���[taT��bX��WG ��rn��<�ِmd���u�a��b<�C,�#��s��U;4��:�E����V��&|6�łZ��0yI�[	ϱ�f;[���x(�i��/RHa&Ŭ����r�� 1Eg�N>Z8\��^K6�h��(Z+�<Vo�eo0C��:�4�*��2�}/A;T�c*��M�H����Ԓ����iz�2���fVů\�Y
 ����6?L���x��y�o��`�c����������'|F��ΥT�tT۳�͕��v����jht��g��倉r˲����\n0�8�:䩒=]' >ԈDH*"1�gB�� o� c ����D����>X�\m+Y�����!{��E۪	�}a4����@[�_zβr�`�e�%R�t��6�,f�؋{]�v!O^��I]g�N���9�0a���t���g�5��Ũ�������p��h�����0X���7Qީ5ͲO�Vf����aU_�z���y�Q�^~lQb�!ޡ$�oa5y?K��	�~�_�w #�T�Z���a���! ��p����o� c �I���H���~MDҲ���'��e����9�����3��,�P-��2�|�I�7���*����p������{��#�k4���MÙp���T��������S�=hU곬n�ڤ���[U�&�n�.ZVRѿUJ�b��nw;���f=2@�,R����h���X �ȰZ�@����LM[�� a~���;AS�=hU�B����B����K�}i��v��#K�����Ga$N�
��!��ZB��,�Ӏ(�r_���#���l�1�ԀU�,f1P�y�VH��T�<�^~���QD���>��Y����h4c�d5�͐�a����g�cЉ�M�_2t�֟�Y�����Y'b�'=�(� h�H�-��{�^�X�;٬sf.��S�	�D��R��	π2�����Vc2�����Vc2�����Vc�m7���e���zTv��d=�U��ƽ]�S'4��g: k��2�����Vc2�����Vc2�����Vc2km� V
i�T>\��&�'D�,������U����r��<Н=.��E�t�	-�Nb�!ޡ$�o����0�9=uS�4q�
t�DY��b�%
Q�[I�ڂ������ iI.s��4w��w������?�z����j�*�����:�|e|p�`5�F$���ɡgJ�w]ᕇ�H<J�B@�+�\���͠�z:n�\#z�`�>���9`�p�0�c��Q"\��M���kzPST��*�ۛ����[98z��"�����P��G���x��+�<����s �s���&�F6�u
�7_Ћ7� ǆQ�z�וyƝ!z.#C�.Y���ݻ �LfE��K�F�L/�x3�TjV�9�3OZ��[/ ��,���Xs ��s�f������˱C�V���p.Eyz��eU�k�7 �TW>PL�t�Aci�n30�A�zc�G@�����Z����)�1�ԠֱTU� iI.s����lp�����2x^����=��klʟ���Q��:'�T�SY]�:�̑�z���]�/)������E�k!�_S1�����o�>�5�Ǜ��k����>�lIorǟD�uiM���	�fmt����]$�﹈�i�~�Ԣ��D{5���U�L�#_��,Vit�-kݔ�yN{-v\L��"��#nS#y����m�(�����p߷Td��#���~$�q����!��ZB����=�+K�������үf�D r�f��h�3(~s)tK�h�RZ9�Y`�ِ{o�7���B�=�7�V���үf�D=�
�a�� D��ﺣ�i��¹ ^��y}$�)`� ��qQ��R��-���fx�Z�0�ԋ�Ƭ�����D�� >r�Z	�P(��$m�&�i�д �rH:FH�O�T�ɲch�b�����#~�@�^l�Y]���p�ݒ��\���l!��'��K��8�0:�L�G�Y#��yl7c9S��D�j���r���4��$���K@�D��;% ���Wy�N��ѱ�+��b��VAoh�!5M�YYroE-�J�龂��K#�u)ɾ��`���i���*ú��-˄�_-��U�4��e���D��ܒ7}p��a~��חo���ܧ�&ٔ°�k�`���D1e>���q�u����,:g�BKV��qO5�j�*Qtu�H��|���f��[����/Բ>�kB	Q>�V	΄,�H'u$�Z0����p�)�����^ڎ�3ŮH�`�|��K�zⲺŜ2m��iH�W�J	����]���y��tq���=<�HI��U�4��ej�3�����Z�N�>�5���Ɔ&"��U qKj;M�̧��v�����e�����9�uTm,0���_�I��O�5s�]�v��8�C1�OԐ����חo���zsلx1=��[|��w��%�8)���r}�Wq�OU險"Yav����yЪx�պ go?�N7�� W3F�������q��1�G�Qc�k]m���yY�A1���X��֑xGV�_��xl�}r�HDʞ�sB�_>"E�K^~��TCZL�d��K�^ ¤+�9-�i"'���Xw�j�7��<�0��J`�|��K�zJ_�xd��j٥P5���rs�i���s+�G��L��>����g���ޔ���Qv����W�Ljѧ4�׿WQ�GG<z��f���$�Xw�xo�A�¦P�.�!�o���m�&�2PZ���vOÉ`_��m��c\Ef�>�77�qO!����C�/7���L>Q;�im���M:��2�n�ڤ���[U�&�nШ��&Q;���@%:���D{5���U�L�#_��,Vit�-kݔ�yN{-v\L��"��#nS#y����m�(�����p߷Td��#���~$�q����!��ZB����=�+K�������үf�D r�f��h�3(~s)tKD�m	$��WQ����VR6�.�3��P��B"�u�߅'O�%��<��2��!;��s\ڽ����	T�|�lSԃ�����d���"���
wh���X �t���(�x�_S1�ޘ��]��Kо�Kj�_���|�/� ��~�̿�:;��ަ�߸
;.�x��Og?6�������O05 S�s�l��&���'b�'=�(#�/�X�?���&�h��(�v��#K��pJ�V�X���7Qީ5ͲO�Vf����aU_�z����6��P8� �+s�ɔ�DY|5-��Y���}E��tteMh��v0<¡�ʱ��VM�d�ꂕ0.p/��sH�}ˮіs�����������,hg~W#_pCeu��|̾?��CG&3�-��_��iz�2����}�u���X�!*�s����v`� Y��(�y�)�E^i�u���L���
�V(k�עi�g���h���R���G)6��	�YI܁��Sq�#�-��'��O�c��M]l]�F7�Gh�C��Nj	
�迿��!�y3�/q�����;�
�{�4'��Xo�m,��"';�#��A	��e��Ż&3�-��_�Zl�<��?�d���&�D�;E��#�g��d�@���;�
�{�4'��Xo�,@� S�J �+s�ɔ��]����ڙ�k����ˇ�������r�G���Vem.�g��A�i�YW�S7�.����~j^�q�����f-(͕2�e(h0]�P��T��zw�\�ڧZ��7*M��J�<>�fpx���:�5Ӡ�q	�۝��&3�-��_��iz�2�nU>���g=��"�ԭd��g���V��&|6�łZ��0yI�[	ϱϲ�ΥT�tT۳�͕���w�����x0�Y��]&(K�Tl�;���f�����q9+t�}Ż�&ǥ��G^��w�&��E������;�
�{�4'��XoN���&��'��P��+BY��9�45��\1��jHM¸�k��CE]�٩��"�@�17ա1�\3�#j<��#����T���{�غŋ��6?L���x��y�o������w_	c��?:(?i˸3�J�
�M�'٥��gVا�˓#��͙�Og?6��m��"���@��b_їE����ݾ-/���b練��Og?6��z��"������@�a�ʢ�#vޖ�C�!��G�*s�D��	�LÉ7�tf�3�%Uo��� ��7CF��ܐ�}�S��/:+�e6j�"Hs<�?j=Ծ����dڐPSn��7i n�]|Y	@
�KS�'|�:w�`�w^���\�}+���Ã�&5�/hshf(�`�X�G[�{�[��/��5�P3 C��ґ�y�x��SrȎ�0h�5eו&��E������;�
�{�4'��XoN���&��'��P��+BY��9�:�d�~&3�-��_��iz�2�nU>���g=��"�ԭd��g���V��&|6�łZ��0yI�[	ϱϲ�ΥT�tT۳�͕���w�����x0�Y��]&(K�Tl�;���f�����q9+t�}Ż�&ǥ��G^��w�&��E������;�
�{�4'��XoN���&��'��P��+BY��9�:�d�~&3�-��_��iz�2�nU>���g=��"�ԭd��g��[;T�!'ؔsy1�n��뾦��"L?��٠����w_	c��?:(?i˸3�J�
�MɂMv!���x�5ߧE4��H��L�}wy�㱏>1�gB�� o� c ����D��n��2��F�0�ε�ތ�T>\��&�����bا*�W�Ǹ!2�͞nOY�c���ta���Om��g��%��&��p�h��в��������eo�0�ܷ��Vem.���9������J��mE0�gǞ��D�r�c��ْl��]�Bcl�/ ǻ��w����Weu��<��E�u���t��>��aM0��x9@xi�n��\ؤ�z;�R����o�a���ݲs���+�%��}����Ғ: ³s�Q;�m���y3�/q���d6ʶ�	G
=�HP�&`&����MԲ���L��S-��f�rE�X�e�!��ZB�&5�/hz��"�����P��G���� �[T�-�"E�Sq�#�-��� œ�ĘK�+���w�����)O��&�h��(�����9�;{�����ml��Ô�R�Q��=f׿����q�>�Yť`�MϦ��pCeu��|̾?��CG&3�-��_؀(�2�x@�����t��y�|�q���~�"����7Xa0~���;A���g�R�"i�g���h���R���ɢ���ڠ�Q;�m��j"^�����ϖ [@wPcIn-Hzn�!��ZBU��<7�9�֝��{�EG ��Z�!3�jQ�V�W�<l+�@EWMT�R� ��O+�>(�g�h���X �&Nm3l�����=�\[Lq.�)�l�dtO��F'ot#�r��8ߍ��{:Q���GljJ�����v·��~U�I�cE��/^�À<MN2��΢�~v� 1�����=��s��&�h��(�5�P3 C��ґ�y�x�Q��C�������$s7A�k�6��� ������>{�w���q�� bާ�kU��r#�-m�f�����I A6˃rGH��*oIt�����*d��ʦ�z6K|�@;��o`��G��]_$A�õ���&5�/h�t���(�x��V���;Z�����.�@��>�̑�z���]�/)��߽����s9EJ�������O��K�fpx�ɥ�W	�s��_��s�֙B���y3�3��(�Y�/(K�Tl�;���f�����U�ӿt�pd����Y��'��e����9����\(iz�<\1k4�݄e�?�d���&��ܱ���wm*��[�!�u�����'Z�[]�g4{��s^��I���=;�������_��s�֙B���y3�3��(�Y�/(K�Tl�;���f�����U�ӿt�pd����Y��'��e����9����=�D����;��|BW6�ƾ��V��&|6��C�jW�8��!$��ck�Bɉ���o{�[��/��5�P3 C������9�<��&�Rȧ� %�?�\�`Z����<Z.َ���'S�c=k�Rm���5���٠������$s7A�k�6��I�ߋ�X��WG ��M�C:4�֊����9����ȶ��Սόѓ�4�LÉ7�tfƧe7��
`����0�E>r���l��˓#��͸t���(�x�_S1�޵�_չ�ŉ���U���Ƨe7��
`����0�E>r���l��5ߧE4��Fi��|�R��G��3Ah	)ޟ��E.t�