// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


module stratixgx_lvds_receiver ( clk0, 
											coreclk, 
											enable0, 
											enable1, 
											datain, 
											dpareset, 
											dpllreset, 
											bitslip, 
											dpalock, 
											dataout,
											devclrn, devpor);

	parameter channel_width = 1;
	parameter use_enable1 = "false";
	parameter enable_dpa = "off";
	parameter enable_fifo = "on";
	parameter dpll_rawperror = "off"; 
	parameter dpll_lockcnt = 1;
	parameter dpll_lockwin = 100;
	parameter lpm_type = "stratixgx_lvds_receiver";

	input clk0;
	input coreclk;
	input enable0;
	input enable1;
	input datain;
	input dpareset;
	input dpllreset;
	input bitslip;
	output dpalock;
	output [channel_width-1:0] dataout;
	input devclrn, devpor;

endmodule
