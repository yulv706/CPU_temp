��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-Ǎ�x�"Ec6G̑�|̍Df�z�g�����#�=�[.>��$^���?�G�P�U��:����E;�i�:��ꄟ��;%�"&����XX�Q_f����N�=1��1��ʀd3��ş���L:�%����:}�8�(�2JF�E�bU��_#`k^D��ń�"&}*	T��(��gjq�=?ل�Q�g��6��ە�q�G@��LF�+,ߩ��A�^����*�^����A�F�7���3�GXS����E@��~���($�J.���
��'p�@��rB�6C�2��G�����#��%&�� ����q��>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z��r9�3�X��-�`V-u9�`�jݭ�F�����K-psܧ6e���Vx�ӣ�3�9����Σ6��u�_����+����U��M��f	����[I����,Y[��FzBR)�5,F�ʦ!�_k�%w�_3#ڸZ鎬����Ǟ��݈�Z��l@+�v�~������]�!��	Ǹ�y85��r>?�W�p��HM�e��`y���9��
)���l�F~�h_3#ڸZ鎬�������(���}/A;T�c�owђN�~R�wX�աzZru.��'���'X��6�vg;Je'���Xw��%�r �&M��y��Iۊ��8���K(��z�j�;9�e����E�$��1v=��`x�~�I+�?T�]D�9�ϑ��[�֖�9x��i��&��TD�Y�J7��e<�1��bÌ�s��X�e���V!���IÙ=�H�^�p"ORmHX���׫�J��q{�f��a�:&�>��s����ӓ��^hq��:�}0�st&���\�v��Q���K�c���%��a�����*�����Ѣ�{l�f|�ό���.ӗ�!����jT%q�#�<��z��}�Q2�+�Y�slxSwP6��B5x�S<��z��}�Q2�+�Y�- 
�@
���C�����7G#+���[H��Q�$�k\_x���� ���J���_����A�2��G�
��吃1�ﻋ-���C�M��N��[XJ[]WQM-���G�yQ��Z鎬�������(���}/A;T�c�owђN�~R�wX�Շ��uj�*��MN����!I/�������A��X�@�5��6�l��s�����[� y�~��ż3���F����T�O�H'�J�����=<�HI����>�W�_=��0���̏�u�=Cm�v4��61��7a	�����Y�
ɸ�oƴd��t�'��9ܛ�	���V[�+
�l掝�K\m��U}�	|^�׽R�s�DH}�_z�9�E�\����8�i�`!31u��9x��i��&��TD��E-%Jn��ɧ���7�)a���%}D�����!��g�-��\��OA�=�~�]��d�Y��o�6�֟�Zl��F�������WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zl��Ͳ�8�3���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂��(%�9>��!E)ėתJ�#�P���(V�0r�����K�9y^6gVW���%@�~� ���I�����+����>�G0�Y���ծǦ�3y
�*����zEK#�E��Ǵk�?H�$�IX[��O2<������ #M�)��u��`�|�&�#�E�d��������y��Ld_���1[���K��&�|�G�2I�wp(��C�712��}ǞK=<^��`Y�F�����I��#��
Mcu�T�M�ڤ [�f!�)�X�j(�� ����n�
_��q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r$����Gd"��U"�̩��k&Q��8�'��j^ҩ#��u1B�c��4`�64�]��Dq]\�����@	Q��[�Fc�k��˚����Z�ײ��Ti����E�$��1v=��`xx��?�&�ْl��]�B/��v
���3ľ�Yx�<,����|#^�Vn�����'MB�I:׷�Fy�XZ@poEE���%����BC?T�<o�nïi�� T[��m��U}�	�(��Q|3�� �����Y~��`�J�2�G�Mlˊ�jJ#�}�����О.�6	O�d^�)�KD(����m�D�c��Q� ���8�%j���V�2�.��=")r��awf��!��ZB���'�u�O�4���u�P�HS|����9���H M��� �\&A(`#+@�@N�%:/�y���
��吃1h���R�ް'���,����%`�U�E�#V�e���锴�;��|B�I��p1o����n�'���,�b�oB|�,�*}4��yή[*%��J{�+�M�( �(�����!.�&˹���~����MA�q�m�,&H�[&-nD�P�E6�Εq�8�:6�m9�M-���G-_6�j@��(KǨ�X��WG ����h	3mi
�,wLnƲU�k�
̲�ΥT�tx(�i��/R��u���NXhA�"���߸��S�ȌsĈ4)'ƲU�k�
�^6N���&��TD�s7�m�[� �3Ah	)ޟ����9���~�h�!�e/����&��e��9�n�RO�^l������4�Ʈ+ˀa�2��Ү�a4�B��ٴ�s�1c��t�R_�f֜��9H�Y���2�x��:*�N�e� p;��w�����]qs�)�*6=�z��f��@|QH˩+`:�l�ޜfb`\�����sB�ǭ����ob	ZH +l�utO��1�Z���t�K�"i����
��+�#G�ۄ��O���azhݪm����Y�{'%s#K�v]|n�aC�h�>�3�nv���|���!vGmZX�t�%&�� ����q��>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z�|=8�E<��FzBR)�5,F�ʦ!f�ӊ[�k��!n}y���q���U�^�n��Uh��w%e���{l�f|�ό���.�cIn-Hznk��HDL|R��{l�f|�ό���.ӡzZru.���/I���g��TD���9�,�w� �:&�sSs�Ǆo}|��XH�����,>$<�խ5�P��9x��i��&��TD���W�5�{ZN >����XM�{,<!W��=Y��_Q2�+�YɢX�B���yή[*%��Jg�)
�R��d�٣��.���ᣓ�T�?�~VOږ�A$�P�U>R~�|L�0z�ͣ��m�twݕ�w[�KX��ik9�$ C��/}>5��0�x��y�o��4M̍���o�γ�hI/��\]�3�� �f��Q�����OOfM�n��x{^4��*m�9�d�L�o�{�R�_����xQ�n
V~$5�j��1Oҏk�� ���ɛ�?ө��h	3mi
0z�ͣ��mbr����Hp9����˓#���5�j��1Oҏk�� ���x�ԉ�>��h	3mi
0z�ͣ��m0@�d>4ޤ�Hp9���5ߧE4�훬�pP��K:+>z����ϰ�ҷ�	 �5�X��WG �����ž����[f�@Y�Mv!���x�����X�@��~�1*su�y�\��կ�ɛ�?өT۳�͕�����ž����[f�@Y'٥��gV������X�@��~�1*su�y�\�����x�ԉ�>x(�i��/R#k�˟ܒ�o|k�Lb��˓#���p��U��	�<?��%��Ǉ�y�ݾ-/���b練�5ߧE4��������*��7�G���L�Y&�l�5����- 
�@
�_�-oH;�A�߹6X�C>�#=��ܐ�}�6߳v�F���'��*�!N�'�y�G