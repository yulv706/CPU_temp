��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-?H)t� �hz2��ƿ� �lJE�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hp���Ť�Mn��X)r����#�L������5N�1 T�V	�tL��	�{�Κ$M�C7y���v6޿���kq����Eֿ�o0��ܧe���5�/���ׇӭ��!�`�(i3[�"5�QJǊö��_��i@�{ۧe[ғr�,�Ōt�}Uٱ�g����.E�^~_|�����{j�G:� ��'��iI+w,A��4�M\���Z ��a�O>*���
��#kz��GN�P�0v���uP!ߌ���^����Wړ��]b�=#;6�#t����nB3�+{Cz��3�<A��d�]��<��&�gG��Hc�e$���=�(v
���O>E$I������T���Q���!i��ӯ�0���&�:�u0&����x2�Zy����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�jM�1}2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!����j.�n�Ax��PR@?�Q|33�����rqn���wѪ	/g�%�W��{�RX�>w�P���u0�������k�V�99^�)�S��uC|Q�����9�ih\���6�oX��s�At�Ӡ�-������u�=�xs�1����";1�(�����]a�{��ۊ�d�k�`�?��<�� ��o�}a�Còz�;^�ru��e��_$߼
�d�YiUbiX>�"��g��3�G��/8'��ި]M�}xf���T��Mߟy�����n��1��\�p��/L�M��Y�Ҁ����r��{��>ڑ/8'�odgƚ�| �����q��5k�^�78���N��ov�Op����	�Y8�>����;% ���W~�_Y�1�����q[��\�jf)�bdZ0o�v�v���O��q�M�4��{i�etWj%h�W�8������8ٓ�j!�`�(i3p]G��>���<�}��x~QTߨ�O3��\�'�y'��BS�z�5&n��ū��@�k�!�`�(i3!�`�(i3!�`�(i3}[x��8��`��Ć?6�!s}6,e �ǟ=EZئ;z&����+�E�r{����JDn ��a�K�.:gdW(o%�)���;t|������D"�~����p�4���='߰����`H��b/3j!�`�(i3!�`�(i3�F{/���!3~�(Z��GmO��%��}�.����M���5^s1@�&'iKb�آ[�~,ΗG\�ʢ�X�=1�����
�^��j"��Q�]f�p����=Qsz����Iv�.�GzEc.������������X�k=o���Fz�!�`�(i3!�`�(i3IB�]�!P���b6p!!v*!���&fB�@��X*,l��d���F6���ׇӭ��!�`�(i3!�`�(i3 lF�Z��f}�y�F�&��S߭;�(6��3{��|o	���=l"�,�>E��&�3�y�2��J�J�T�S1(_�'�&r�~,ptQ��k$Vʴ8X�S����TXP�e�g]�H��֟B��Ўek'`�j�13*�á)ˎ	��[�!%&oA�\ֆ�
'��(�<��
Aʎ^g!�`�(i3!�`�(i3!�`�(i3�|j��"C���ޝsn?V��-Q	�	:����lg\ ����EO�{��ϫ��u�o���q�Z��?��: 0[�T#�l�/Zw������{%hPb��͓T�)��z��z
��K�O�n���^���D�*�Z�J�v$��A�f�y'��BSƹ�#�y�w���	B$�@�A�w{6��(�N��K�O�n8�[ �n�
�CQYb!��uፁ�&�$`8�+DO�n�;4L&�y;U�2y��}���[N�)J��7)�c�0:S��}1yYZ��� ����@	�1i�myh�~�*�.i,����j�Ə���&,���9�tOHn����x���I8I�%-4o��Iu���'�#&��
 {�L<��-�|��e���RB����bb��Ə���&,��+���!XwOHn����x���I8I�%-4o��Iu���'�#&_�:q`��� �Z)}�6!ת���ېư���o���o��V�x�O`BpI�ҽb.j����kѶ���� ���X%��m�Z9a\������0;8�y�%$���r���{��6;)ܟaTo0BpI�ҽb.j����#�2�/D<�L�k��\|�M4��*��J�Y��в}��aC�2V�Vׇӭ��!�`�(i3!�`�(i3I����Ǻ'n;�>�rY
�����+O~%��짐~��.d����"���p|��X^䀸~�W߁�nrm؊(�[���~$�B2���m���-��
�8���?�*���\�Ə���&,Ƿ	DTjE,���6��q@�2��>�b!��u�Z1~�g]�u�+��
~J[����30�A�zc�RhoŜn!�`�(i3!�`�(i3!�`�(i3�M��n���<����lpU�:�ƅf��	��������6��q@�2��>�o����|�sg�2�:��~�^=��D�,<�V�QK�}�9���u����Fz�!�`�(i3!�`�(i3؝�4W���+DO�n��t!I����;R���fǥ�c⠵���طYRdZ0o�v�V#��ب'�����{��6;<� ֭m�_���ȃEE��$(��{�$�˽�Lk�`�?��<��t!I������h+�w��4܆��O�2C��OG;�['*�p!!v*!���O�{�
;����"����+H]�����˶���,/Pc��?@W��8�����b2�{������7��U�:�ƅf�H��������6�����+��w-���f*���׎o�|��Y�� �k��^��Xz�Ȗ��W�{N������~چ�sֱ"MT}���o�׎o�|��Y�� �k��^��Xz�(��¦�L\�kg�Ť����� E��5�O�U���.b!��u�w���v.���A�I�z�9w+�!J�0©	]�,�\DW.ɧ/H>y7�J�]f7\��1�T�g��������G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcn��^��N�oߛN�N�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hF^����i�̨���qh�'aba�	���
��?��n;�|-�Z��2S ���k��m���$[΁�a�n��Vk��w/&g�-ΘBdN�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��f����om2�����iҢ��V�x��%�a��i�9�J��$b6�]ʆ�In��t@���z������)����")�^�3��8r�Wk�ǻow��R�nI�GI$��ǂcY�~遅��'�:��'n�^0o��S��S�Ib���ό���.ӥóM�˄NQ��臿5"c'��ɿ��3P�d�8!��vp�P}��O���w2T��b�T��xd�Y�I�;\h!E��c�G�*ZkS0��nB�+������]��)`���"��y�LN��K��g����R�<�W�C%c�����<�W�C%����_Wr��;���EWr�L{1��ox ������ �i7�sp>{=J���.��W�}�"�,�>E����\�vūx`��:��g�0�u�L{1��oxr�O΅��C?�D�s�R�"0��<��	��������JF!՟Ր��M�aW��Σ�?��<��z�"�~��S�
/P��Ѷ����A5wr�4�Vgn`��p���n�O�V�N�s
l���u���NX@��^��>��}� ���O%��y�䃶&f�����SVc�5ߧE4��?"����a�m���q�l;1�]�I�rT�8#�>-��;��S������yq]C
R��T
�N�oߛN�N�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hF^����i�̨���qh�'aba�	���
��?��n;�|-�Z��2S ���k��m���$[΁�a�n��Vk��w/&g�-ΘBdN�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��f����om2�n�h޶�\�Ji��'�o��Q$������aU��D�	a���(�E��!�`�(i3l0��F��j���^B_�(ba�7�X��)z�s�!�`�(i3%Ah�%4
>��XP��Ȱ�^�7^/�AJy���l�f�nϵ ���3�ҺIÙ=�H�}ʧ8Еb����������gE�,�Q�^�y�zL͊�q��_�0���ӨI��'���Z[A�E����F�'n�^0oL��pN�5����`K�x��R͖"�,�>E����\�vŻA�1�#`�͌4s+�ny���A�!3v!�`�(i3JHn��z� �&�^`(���%�a�N�+��#�!�`�(i3�b9���6,� k\\1�*_��hc�ʹ���`!�`�(i3l0��F��j���^B_�||�?�5���J��xi��͆'�X%Ah�%4
>��XP��ȵ�d��w����y{¦�$]\� ���3�ҺIÙ=�H�uoglR���c&;�p� ���S�Q�^�y�zL͊�q�� �-8���I��'�	�ų_��E����F�'n�^0o%|�J�0�5����`K��q��"�,�>E����\�v�Qq
˟6͌4s+�ny��9� W0�!�`�(i3JHn��z�k��%��6i��%�a�x�+Vv��2!�`�(i3�b9���
Ay�9�6>1�*_��h���Q��~��
c�[��ƣD��T�����NI�����m�2�Z,qC͌4s+�nycfl��6t�$X4P�JHn��z�S@�z�R3��%�a������?6�9������7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?�ɺdX�-�B�85���%�a������?6E�C�Έ��7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?�ɺdX��<�-���#�p������p:�2],˶�9�c	o'E!��s�Zu�EPD]�I���2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u�m�\��q�Z˻r������U�r�}��}����ހmu�m����y^�k���%H�$N�oߛN�cL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��D���X=��f��i��зq8�ЈxKʜ�#xI+r�� 0�D�A��t��D)��i�d��`m�¨3��%�$�������\O�a�|�6����&��DErwⳘ=�C. ��f?��s^�xct��_Tҥ!�V��NR0�����O�,�WNT�N D|�5N��VA}�v�a'����\�Z��'�Wa�L��ʻR0�˧���.�E����Fr<���\�g�-ΘBdcL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U��k�t���L53�����)-}�vPt�>xA�ꓩ�l;��!I/�������A��1��+�W��J�ݨg4$ _o����OI��@���:��F�b��@�zL͊�q��c�sYIJ8��OI��@�n���������Wq{�f��a��{oS�=wK��7�&d&(C�#�7#^�Vn�^ֻ����XP��Ȇ<�qp^S��j.Z��$�sӢ�]3�����c��(r$����G���'aOދK-\��$-��Ǡ٥L����e]�u�����!�M�T���ݏ��A�!�`�(i3���+�J�������"�,�>E��W��Ґ�YjZ�p��Z����r;��*!�`�(i3"�,�>E����\�v�!�`�(i3Sn<Z�)K|K�@�����!�+�!�`�(i3%Ah�%4
>��f���T,�;C@����%?!m�Az�F��O�4p���eq��VZ�0�s�b<�B�_���X�KM�����7������
�]qE�&���W����Q�^�y�����9�!�`�(i3���3�b���-the��戉Z�T!�`�(i37s�9���o��S8����J� �j��h@S�@�]_LO!�`�(i3JHn��z��x�f7﹏�1β��h����0���,�W�B�޹B$~s%��@�:�����xwƄ�{Ƨ\-TX�Rj�+s�!���r��*y�xDp��T�/i�M���"�,�>E����\�v�!�`�(i3y�Er�)=�ᏅN~z��9�{�G�K*V׹ږ��_��f���T,�;C@����P@zQX�76�$t8[��5��FX9�p�x^/8�D�n�ؒ1ECWI�R��R��=���b>���F9M؛��&�}�(�dW�,��(�a�肢�{l�f|�ό���.ӟ
�r��	G$��R�lD<��z��}�Q2�+�Yə~�yD݃��r��DB�����I�b}Ω:���V�(^��<��z��}�Q2�+�Y�7
�4�.�E����F�ҋX����|P�������A�=�8bH���L��B�;#5d���7Ê7�E�4'���Xw/���:;aR[�T�.�W���1�}�ױ��(@�E����F�ҋX����|P�������A�=�8bH���L��B��)�ޭ-�7Ê7�E�4'���Xw/���:;aR[�T�.�W���1��)$磨'jU-j�`�ҋX����|P�������A�=�8bH��Ę媌�+�<1(f}ظ{����$ <��HT� \r���㯄�����
L'���Xw��RN�-#�ьb2up,zk�g��[��v�$ƪ;���Q��/(A=�kX�*1�e38����2�9)�����m��T��J<�]qE�&�owђN�~R�wX�յ�8�,wO۳�yz�<��z��}�0z�cUL� ���Q�'e����u*w�A	'���k(�պ6<��z��}�0z�cUL� ���Q�'e����-��\4vߖ%��mz%���=a\�&'UR�q������3���R����o秾�!a�v�����w:ꮆ@IE�U��@�ڗe'a�v�����*� ���@IE�U��@�ڗe'����h+������E��@IE�U��@�ڗe'��;R����H���i�Ox�j�d�ƥ4�,�:�'t��t�W�lT[�HF x>H�|�Wǖg3ȓ8���/�A���0v7���V�x�O`�����
L'���Xw�j�7���rcJ]�0ݫ���Uh1�gؘC���t\>��fm��]2�y�Z鎬����)��e���Rf?����]2�y�Z鎬����)��e���= �J4��]2�y�Z鎬����L�`u�K�˱�Ui��Q�x��8�,wO��ٷ���TD��-�`��8�4�%��mz%���=a\�9�K�v`0���'=��"B��$I��w��,��xc�l��m
��5�(�����:x�V?W�)�ޭ-����
L'���Xw/���:;aR[�T�.�W���1���~������yf��?N/7G#+������z����A�b�*܋���ԓ�Dd�<�,E9|.���%�S��v���?�R����o秾�!rF)���X�3c/��!ő!XF3�@IE�U��@�ڗe'rF)���X�3c/��!�:GV��d@@IE�U��@�ڗe'rF)���X�3c/��!P;��	�@IE�U��@�ڗe'rF)���X�3c/��!4V(�x@IE�U��@�ڗe'rF)���X�3c/��!з���jf@IE�U��@�ڗe'rF)���X�3c/��!�f���l @IE�U��@�ڗe'rF)���X�3c/��!�Q��Y��@IE�U��@�ڗe'rF)���X�3c/��!��8�ۦ@IE�U��@�ڗe'rF)���X�3c/��!��A Ly�@IE�U��@�ڗe'rF)���X�3c/��!k�O�`c @IE�U��@�ڗe'rF)���X�3c/��!����4��8@IE�U��@�ڗe'rF)���X�3c/��!.�0�;l@IE�U��@�ڗe'rF)���X�3c/��!'��t#~t@IE�U��@�ڗe'rF)���X�3c/��!򊫖��@IE�U��@�ڗe'rF)���X�3c/��!��];p��@IE�U��@�ڗe'rF)���X�3c/��!���L���@IE�U��*�QN��� ]���f��v�鳔�Ċ��8���K(��z�j�;9�e��L53���Z<�~�q��]3�����c��(r�CRQ���E�+d�ίp��V�����Y����딼�\�v���T�©�#��l�َ2c�'z͌4s+�ny�X��{��ܛ�	�����^�%k IÙ=�Ho?Y���	3�Ð�9�X�e�B���<����ą~c�PƐt
����������\�v���T�©@���U@���:��F�����XuY*"�nw��F�dZ0o�v��CRQ���Eu<�.��	�L�t0{�A����8V�l0��F��j.��h��u>1�*_��h��Ӯw!)��&�t5C�,���m�b9������U.6����sd�Hc�.2��w�k#�J����͌4s+�ny\D}��^�y�����"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s�6F���y�8� �w� G�"�|� }�Ri.����l���r{����JDn ��aů�x� ���rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'��KD����w�Ve�U�ԝ5�͌4s+�ny7\�%Lţ}���u=|�z�)�]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s���A0�>�8� �w� G�"�|� }�Ri.����l���R�0�;"��9�{���|hY���rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'��QV&�f�w�Ve�U�ԝ5�͌4s+�ny�y��P�p�V��O"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��{_8�Y���˂lq��r'��i�B�J@�l�s[�5����`K��D�	a���Ӯw!\�8䮨��ekW���I|JHn��z��ea���4p���eqd���w&�r��VYW\�����[!�`�(i3%Ah�%4
>��XP����~��84Z�Ћ�l�TE�խ������S�0ů�x� ���rs�i�Vw�C�-��0#�tC%Q,!�;��
r7��(*h�Qf�kCH`=Th=mP��T�͌4s+�ny\D}��^��ٙ�D�s^E��S�Z鎬�������(���E�̱!\Z>�
6������+$��g��U-�e�v�W�G�[�^�������-the ���mh.�]����GC.�|���~��H��efm�0z�cUL���a��<mDrW�B��"���PB[<b�P�`<����B��٥P5���rs�i�H���N��C�X<� ���B��8�R�Z_.΄x�g��	��S8��UV��\Ƴ�r��Gh�Qf�\l{�"7�sa�vݝh�c�A�L'�1�d��{�ʬ�缆�YW)��͌4s+�ny �Ǧ�_@f���_t��R��XP���x���: �&�(E�{�ʬ�缆P �8�-�US�����U[�[B��$�����˔b�7D�EI����I�O��\�v�d�jFB��]͌4s+�ny]"Jׅ����d��.%Ah�%4
>��XP��Ȱ�^�7^/��1������p�V��O"�,�>E����\�v�VNub��pzl��a�Ʀ�|þM��a��zr,/'���Xw�j�7��r��&D�:f��:F�X?�g��U-�e�^.�@���e��0�U+�qbp@���K�Q�f�;�>)ʁ���f��Y�{'%sgeߪ�{ ^�x~�(vi�t�c,�q�T�\ ��-3zYIިuIF��^~�$�x�Wt!�`�(i3���+�J��Y�{'%s���䒼�7��Hn#���T�\ �͘�f��p�b�z'hۉ)���	4ˣF�n�5��cz^8������зq8�Ј'���Xw��fi~�'K�2��J���"�!ɺy���B���Ȇb�L���g�"�,�>E���]�!��	Ǹ�y85����@�`�8�Wǖg3ȓ8���/���fi~�'K�2��JHm����v�V�Nt�s$]�6����ޤg��c�n�5��cĭ#�?UM�!�`�(i3зq8�Ј'���Xw�j�7����o_��ü~���U��g��U-�e��)���UM`���R.OƋ.]$�t_-Z��T�\ ����Hq���F x>H�|�j���Iq��w�Ve�!8���\/Üy�a
�:�,�!��qƸ "g��z�WCp}��~Ϙ�g����P"X����G�"�|����.N����=��Ʒ����V�3��yɶ7s�9���o��S8����iY��"w�z��C���g��U-�e��)���UM`���R.���b\�#@[�I��Bg����P�ߪ��w��m�C�7���s��R��һY~����j��n�t�q�ٲ��+�J��Y�{'%sAX���	q���b\�#�y�Ya�I��g��U-�e��)���UM`���R.���b\�#�y�Ya�I��g��U-�e%uX���4N�|��Z�<kx8냞�!�`�(i3��Q]� _Fr�����WF!a�ޅNA��6D���K�Q�o{��:��(�[�*��Q]� _�rs�i��O3JT�!I�T�\ �͘�f��p�b�z'hۉ)���	4ˣF\d�RI��������yبw�ሑa7s�9���o7�B�J���o{��:�N�#�@j��{�`��Ҝye��B�o�\q�߈q	���S�[N��t�$Z���>�ߜ�J����^�_�J*�(��Z鎬������D��찔q_�pk����2%g�#0~��}�� л��@(�Ϯ(����%��yBD~"[
W���VYLl*w�{	�C�9Jn�+��Q]� _Fr���������0�@�U_� ��*ߵB`���!�`�(i3�!��@y��=�-Ǻ�:Nɲ`wl�����`�Ǔ3zӲ݌���������j��-�n`5�fK�Q2�+�Y�E�!Up-i�Cߋp{T���[�2ٛ�X�/R��:2QYeƈ�c�Z�~E�!Up-i�jK�o[���[�2ٛ�X�/R��:2QYeƈ�c�Z�~5�e`��9d��l����v�}���X�/R��rs�i�H���N��/Üy�a
���"X��[�p C;8;kѶ���� ZkIb!8!�`�(i3�d�٣�����6>�����ev.������f��gy:h+i
Z鎬����Ĺ#{��a'�<� \�Q�w���*��_?�v���Q]� _�:2QYeƈ�c�Z�~ݓ��E�I�Q�Тd�!�`�(i3�d�٣���,�JL���+ޡ)Ծ�/�n�*���?�#�6�fȯ�?
YT'���Xw�����C��'��/��࠮R:������V�6IWJE�r���秹��ч����=ў@'���Xwd�n]N�^ �7�}3��|�b�@a(􆿳���Qs��������=�8;�(�[�*!�`�(i3Ww�[h�q��!���\���Ȑ�'t��t�W�؏ 4�+�{_8�Y��M��)=໺(ӈ���x|}�|0�(�Y�MM��5��g�g�(�[�**�k�����\F�^�	E��߅�'e���婣	���U�dN�<@Iv�H�_��Q��b�z'hۉ)��!��|"/3�+��m\ƪ;���Q�0�=s�����[q�2�ߣ/s����.Y�[&���,�v����z��ˇ�h��ܙ�[-<�+�my$�N��YͲ�pzl��a��Ǯr!�`�(i3!�`�(i3�n`5�fK�Q2�+�Y��׎o�|���Y����!�`�(i3!�`�(i3�d�٣�����6>��i�X��*Z�!�`�(i3!�`�(i3�E����FZ鎬����Y�V��#qFL}��!�`�(i3!�`�(i3���+�J���q���U�pzl��a���gE��҂ϱ��[��Q�#<4^��n`5�fK�Q2�+�Y�kѶ���� k���3�F�-XX!i!�`�(i3�d�٣�����6>����9וP�;xB�_/�1!u7}:�E����FZ鎬����Y�V��#q胬<ċIX3�A���\�J2)V���+�J���q���U�pzl��a���gE��ҩ���;//M7$����n`5�fK�Q2�+�Y�kѶ���� k���3o=�<*��e���b��d�٣�����6>����9וP�;xB�_/]k�WM��q�E����FZ鎬����Y�V��#q�?�B��{k���3�z�Q�q���+�J���q���U�pzl��a�-{�*�;�Eo��K��]�q��n`5�fK�Q2�+�Y��׎o�|�8����|�M��5�!�`�(i3�d�٣�����6>��P��r��c� v?b���7;�Eo��K.�wK��� Z鎬����Y�V��#q{��>]#���)y(�O|�M��5����+�J���q���U�pzl��a�����;kn�P��l|�M��5��n`5�fK�Q2�+�Y�K=J��(��I(ީ���a41h���������d�٣���Ni�4�ڼ�t%>^��?�y��hL5ӥ����c^����
<ڑN���2�A��1��R�9*�eaA�|j?�d���&���>E��*�(��z�¿-ǂ,yߊ��b,�a������)�}�����T��.��W����t�.�!�8�}�\���;A<�SNp>�3������"h���ƅ5����5�`��N�W'�o����f7����e��x����#E`D���$G�	P��?[@S�CZ�~۵�q�#�p�	;�0�e�n�xdɨu �䆡X�dr�jf'��H������V���
���F:_ʣX`��_/��IC:GMG�2�3�A�E'����>E��*	Z�~(jm�7jl�N�Ar�/=�N�}���X	j�w~jiǎ[��S��_�:�R��h�4�b"����gE���Y(��	Q��H/!�Sy�+�z�}�-�%Q�a�4f�+�Z�{�b7�-�4T����	��,��<����r�k�,��~��U?'�����ٴ��{�G��ͫ������:[ۚܖ��`�[�	2�GF�&���#VW�GaAO'��7wT�,���P�&`bH$��>��L��$�I��i�j~>�Q.Ss�@�������-R�X��%�VB�=����R��(7�
��o��N⃟g��|"u8��d�w(�`��l4���/A� e8�~��f��Ԡ8�tF���)e���n�`�v�Q��7[32X|��h�ɑuϢ\�S&��)Q�����{1���	m���N����B�c���7zxs�ްs���	m���N����B�!2^D�S	�o�7s�����-���
0yS_,D]8@U���H#��Ɵ���X`.�	����Y�oc!���ٴ��{�G��ͫ������:[ۚܖ��`�fJ�WM�.�A<�SNp>����AnJ��ó)�󼅯|��%6�Y�JDFH��z���8�ϑ��[���D���0�j�J�Ñ=��[1�%n�@��V�����Y����딼�\�vūx`��:�,�qo�,ܛ�	�����^�%k IÙ=�H�]ƭ��&d&(C�#�7#^�Vn�b9���sW��NZ�uw�@.�/wc1��˪Xk"�,�>E��<��z��}�Q2�+�Y��1S�����Y%T��BPS�)37J*u)T{6T'�f�;�>)��U֔�>V	�]�!��	Ǹ�y85�R�m�.wa�Iz#1�<Td��"X��[�A��N��|�+�� VU+I�z�c�5����ݱ�Ʀ�f�������~T�����A���gf׿���$	n��s��ͫ��;���^hq��:0k�y��HzL͊�q���19TH���8�6:�F!�`�(i3l0��F��j�
����uK9��>�������q�}5h�-tQ���͖n!�`�(i3�b9����6�{@$��uw�@.�/wc1$�W��9��I3���S�)37J*uc�A�L'�	�Vh�/�owђN�~R�wX��v~S*��R������5	��]�!���������RP=	P��{l�f|�ό���.�L�2�r�Ĳo  ��]�!��V�,�q^���ȍ�)0f���{l�f|�ό���.�V�|M�������5	��]�!���sC�)�.;�<.��{l�f|�ό���.���S��"B��$I��w��,���|HH9M\��e���S������
�:�e�ӎ�4���S������	�_���X���n�k�r�>?le��pp��]�!����-joG�j��ԁÆ�7G#+�ǟ
��|�6�E�W#��e�0
A����l_�U�x��3����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h�����7�$�G�j/����X�e��}c���G��m\Ӓ�qܛ�	����(:��=�M��0�d�Sd��_�a���n�|Wg�|bVzN7	+`�9
EMܓ���;�e >���l�n�Zl��Ͳ�8�3
�{�-�>��t��ԱͽP�nT�_ɷ�}���y�L*���8�^�.eO��q��S��;�(e)��v��=����'�$��u,��y�"���Չ-d��r�b+��/6!��Ei�gz�����n�|W;"V7��evwJ���&�o�\,9o$aϛ`!�A���
+,I�2Sj�	�$ɜ�\�۟�-?�d���&����{ԕ�h7�{`��������* -��ed.:E������ƄH����[��2����s�ZK5U�㶰wi�G�A����`�+N'����)�!9x�����A��Y纽|ԯ/��m�h@ѐ�ER�)��<|+!N�e[�������C1�у�ӌ���qfb�B�l�2�����^t+����2�\��v�"f$^���\�}�J2)V	^�����v���?���1S���������;q&1f9m�҃kG���!l!�`�(i3W��N���;�������<�K�kσ�a��R�#����[��G��mO.�����R����ć��mRiP���uVw�������`�-<�B<.A���0v7��)�ޭ-�΃$%HJ�#��|�k�HB���15�-�bFd%��I(ީ������	��+?�d���&�Ա��+��i���%Ὠ���0��H22��=�z#����2av����pJ�B�	e�q'�D؉��_�m�����W���9�b�w�䩳J �s���H@�{���]K�I[;;v�W>�.�5�O�O��S�7����eߖG
�<ݬ�K������,����k�*�.�a�n'�,+$\�M����F�V����Z����H�ЫY3EZp��Ĺ� ��p[�ٕ����se�{�z��x� ]
�"ǩ>�)E���Z��v~S*��R�J�a$�Y 	�z��V��2�jE?d�1S���������;q�Y�f�ƥ�d��Ke�ά@�ș�I����~u�B�f��.X���ֻ�����h+��
!O:0��O�W�."��ђo�N����C����N���&U2�S#:�*a��E��]n���G�87�]���`�-<�B<.��U4�i%���;$�{�R�$�V�o=�<*���Nm�}��0����8�D���"��	���Yb�V��	��y ��f"�$�!����L�����©h\���k�9�����/	è��0�	+�����6(���j��h@S�@�]_LO�Ŵ#����#g�k��m�z5�Ւ���Z	L�'�}5� }�	��%���K5U�㶰wh�(R;�����3Y쐅�	|�Gy0E��*����	��۽IM>�������ܪ/���ܸ���$�;�5�sw���J2���;B����ՑK�^��F
f����w	}��tsb�?r	�'3���EK�����
�F���LS�ߛ7�C|�L����5uE�(��*O)�J�1U"��2 9�Q1~����?ON���?�� 5傟������kV�U~�X��9&���=/
��G�~7��|YYp��]��nq/����[΂8�:b|�%���,���D��\��%��	��<�T?N�·�����9ۇ%p� ���3�y��9�<�{Pkt����^�r��3�h�|��4-�Q@_8X��Z1~�g]���f������y	��Bo���+�hi��;	�v�鳔���bL�%s�^�� �	���bl�����7�-m��0����NF>4P��)���=E~���e����
��M+)U�D���ڡ�$��2H��&Y��V�'��С������$}%��oR��ן�/��-ށ� ��*lxi#�3��|��4-�Q�p����i�7-ڍ�mI�ｘA ��
�A�m�`�H_�U������%Ik�cIƼ̰�m���;��u�(�};�1F�]�q:�q���8̈�f�������,�Ȍ���\�H�f"��ɔ!:����kݛ�l�a�t]p��Ү��~�[_.H P��?xA4����2��<E눏����ܪ/���ܸ���$��L��ߨ����f��C�쌓���2�����=S�vʐ̡�&Y��V��� ���)���F��=��'?$���0#��=�\���@���,2���!*�؍�~X��a@=�����Yx��t*�=a{��67�M��(�K!2�7�&���=R��
G=�H�쭽�o����rN�>���t�'%��H��܌z)-t"wdC��_m+ �����*��W�Kb���Z��KD�И|��,2|�Z�F_u�
!O:0���.�Ҭ�^}�]���k���3�F�-XX!i�N���&U2������PG/�W���LU�L���)�lV7�]���6��(�N�3���?�xB�_/1d�H�Zc�{�R�$�Vִ��l�+,@�uU� ��}n�8��D,�K�-)K�'h��Q�C��1Dm@<�9�X3�A���\|u��W�s ��9�Q�Z^ >�@�uU� ��}n�8��D,�o�fy'h���I(ީ���x�tO7����[�����|\���sIN�vvH����k����ɝ\�!2A8�r<����P ��BP�wb�H�Z�^6w��<��D0m�'1{{!LU�L���n�Zm����)0kcj1�kD�t�Sj̆���K�|�'�ȵ�]u(+֢���S,�D�c��Qԟ��
�A��R�j`D�����4m���Wӭ�6@ri��P-{�*�;�Eo��K�p��h׬V�!+���}9��m;�n�i?3�(��'t!���Ci嶨��V����m�=�er߮�Ȗ�%T#�5��gE�����b�ђا�0�)_��c%����lxb�뤆�J�e�C��1(�����d^_�Rꑽ,�I�d�N�1�b�*�4MM��Hi嶨��V����m�=�er߮�Ȗ�%T#�5��gE��Ҁ�M����]��Y;�c%����n������И|��,(�= \	\�M<̜Z���wt��B�A�M�I7g����i嶨��V����m�=�er߮�Ȗ�%T#�5��gE��ҩ���;//��0�)_��c%����yg��c|q!И|��,(�= \	\�/��������Ch@�����y-�c��d��ȵ�]u(+֢���S,�D�c��Qԟ��
�A��R�j`D��R'�u)]�t<���J�?�� w��l�iu��T�U9��
�;�Eo��K�p��h׬V�!+���}9��m;�n��(��H��_�0��R���־�U��sp֟kh�W�f����C;��҇И|��,��N�i��!��z�w��<��D0��8#���#����a�9�;�Eo��K�p��h׬V�Sy����!�`�(i3w?�W�S[И|��,"��7Ch�m�1S���������;q-{�*�;�Eo��K�g&�?�U.;�<.�����^��1uv��e���%�G鉖�;�j[����"��8�O_���`���k���3�˙	e
^�I�*�y����(@CPwn������И|��,"��7Ch�mRiP���uVw�������`�-<�B<.�,�I��
���Ƀ@tl��(Ur|u��W�s�ַ
���iW�\G���J�e�C��Lle�J��0����1�T1���T^���И|��,;�L�����G�Ȧj�v���� έ��F��#�Ц�w�L�������"�$�㔩?'�m�6X���(��ޭo:��gڳM뵨�I6�j4̗��W;��"r뾃	��s�Gq��M�B���޹B$~s`�� �:Ft�EO�{����O�2��a��x))b�K���$73���'���)E������?�d���&��n=:�Ed~z,�	��lx��`�+N�%'ף'���i�7�^��X��=����`�+N'����)�!9x�����c6�c��A>	�x��FR��GN@����x�hn�B�l�2�����^t+������\��vMjm�f����qfb�B�l�2�R"8�{����=���z���X�v�J���C�O��S�7���޴:�Q�� +@����T���!�
���qfb�B�l�2�R"8�{����=���f�H�Γ�^���\�}&�1d��̺Eh�m-6�c�����0�J����<���r�G���6���U6!w����}q����߄1�9F[0�#����X��=����`�+N5|hy	$��EV_�[(����R�?d������?���+y��"nF^�{��s^��I�$nx떖ݏ��A�7���?�!���bJ���WW�+���3��0��A����}�ʩ�Vh�l�G!W�:4'.�Rי��3��0��A����}������T{�o�����'N U����k�*�.�a�n'�|��1�)�S�������Z���b}Ω:���DIMBg�k� �%[V��	��y����}���H@�{�'IK�L�����d�k�;�r1΀�]�n�H���E�K���_[�xT�m�Ht��;��� Ɍ��<�,E9|.���%�S��v���?�R�����&���"����2���r�\{�j��?��A<A۞h�G�!Is��� ���,�qm�c�,�[`�&�뵇�@�;�H���o ���Gƈ2�	�i��#�f�;�>)��-��Zz��캧xӍ.��;�N�cP*{+;����'�SS��[%�lM0�`NR���c�,�[`�v� ݼ��rF)���X�3c/��!�R��:�}�f�;�>)ʷ
�4�� ��R�<lͬ۞h�G�)�|i�l���I�&�`%@�`�4�+KK� ^���PG{��_������
�]DWl$�`�]
���b��Ĳ�������2�����ǈݻ�N�E�Q3�۞h�G���Hz-�O�R�<lͬ۞h�G�U�_�}A ����I�&�`o��Ow;t4?�C<xWY�K��e�Igg�6��@���DZܤ�jM��3�}�v*��;��g���2��<�`�hE��Ez	*HD{۞h�G��~q�e~B���,�qm�c�,�[`�[��myAp��;�H���o4Go�HHm�	�i��#�f�;�>)�,Զ�1�J캧xӍ.�A
��z(��L�(�rY��'�SS��/ل�� `NR���c�,�[`�Gh;ʹ�[�rF)���X�3c/��!� Rƙ7�f�;�>)�-m>c.��{�	�i��#�f�;�>)�:�l���i캧xӍ.�9��7�_�g��T45�y�U��䴃���%��������n��\jɖ�䴃���%�������c�A�L'3!�������p�Ӧ�3q��������<iKT>{�ׄ�=����%�[�:V�J��!�B�b�x��h��B�
f�ndu�Z鎬�������(���^ �7�}3��|�b�@a(􆿳��_����OO�;���EWr��;R�����a{7?7s�9���o��S8��<��Qʵ�]qE�&�owђN�~R�wX�� N��r*��D���6B#����߫UӇ��ɋ� ��X�D
CvK}D$>Zr���~u�F8O*�E3* �s*F x>H�|Ċ9DX��&{H�3)-(�K��LZ�|�b,��"�T6Ͻƪ;���Q�����̅�Ż�&ǥ�̻����.�(�K�t�{O�v�dI���}��;R���~��R_	P��u���NX�?͈b���l�&�Yw_t�'wh���R'cf����(-ЀU�D�� ����ɵ������a6gBa�����0�Lz��q�۵�ԬFi��>��J�Ar��� ��o_��ü~���U�z�"�~��tl��(Ur��뉶�N��i,�	�����;R�����a{7?]�z�g9w�fF�5.]��۪	�}a��[�.K3�$�)�vx���a��e�tf���!���!Qr�g?	��ofob0�۞h�G���w��z�=k�Rm�����Ʀ(c�,�[`�z�����?g�d�)�QX�&�E�K�~V��=E�g�������(ӈ��� �3�c`�k+Q�h'�Ȝxڣ9�$���>��o�����}�bk��=��bݙ��N�g�c�`�B<�q��L.bC��U�gQMf�Ʀ�|þM�I�=X�����r��Ȯ��ߊ�u*w�Arw�&�z<a��N� ��M�W8߸��S�Ȍw܁ZUz��F�Y�ɒ�I���w��T��? �O{	�8�to��h�T��Ƨ�2�juWE;p�̎�)6Op�/rCq|�ْl��]�B}Ю�01�߽K}��׍�������x���y �谝��X�e��~��qRmHX���i�k�Zׇ	� T[��m��U}�	�(��Q|3�@���U@���:��F��:vP|c�PƐt
�G���خ�;1?�[F�sp֟kh��*�T�P!�`�(i3L��S-���g�rz[t-��!������e'��ǩ����M�۞h�G��;v��{�����h:v���r�M8�f�~�/i
�\ ��.rV֡�;�H���oor��	P�ޓ��-�!��Tӧ~�;�H���oor��	P��1��X��WG ������h�v��|��Š݄����Mv!���xԌ��Ǐ�c���w�I�7ݟ=�NM��40N�J0�ʂ�j�Ï��	�Li4"�	����-���S�w҄ھɲo�I�xg�~p!ۓ�x�DUJ�u�q0O�*�]��	He"��Ç�q@/��r �����-���S�w҄��	n����jҵh�f&[�>
�2���fp.͏�����6��,}�,?�|�cc����{s��,�9�{��(%�95�2]y	:���a��d銦�i"�S2G�
 V0�zc�,�[`��Hm�B��j=/x9���G-�#Vl-�	�yH@�
@����=7�}|��	�3�� �f�u�q0O�*L.bC������'>D��O�7C�&Ut�\�����h�v��|��Š݄���'٥��gV�J��Ifq�����ӮvZ=�9��f;[����\�G�����z 7	B>�b��O����~y�
3�V��p����<dh�}3d�jK�o[���[�2ټ�mˊ��դ�Hp9��Ԍ��Ǐ�c���w�I�7ݟ=�NM���x�ԉ�>��˓#���J��Ifq��u�ǏX��=�9��f;[���aS %'`m�6��HHD�u\�!�p����c�Z�~rw�&�z<aSm�6��`4�04�jf�5ߧE4��Fi��|�3;c�<�3�Y��jb��Ck�8'��d+�����C/:"�����j�_��l�؊9�~��Z2��r�a��A�q�̈́���#~��T5u��@���*�n �_�:��ˆ�	�(�����+4��v�W@aKq\v��4�s����>Y@#$Kb�i�t�G�|�by�R�QY�v��|��ź��$�!$Y���@�}Wq�`ASβ�=&��]
���bO��Ӈm�s�F��� �h�gc�>� �_�:�՚^&u�0yf%���G����.��@#$Kb�i�|i�&���	K$�ْl��]�B}Ю�0�`m��';��?2^�9c�,�%Dvˊ�jJ#�}�����О.�*/���~���;A���g�R�"OL�Wr��{�ol�B�IY�5����Ң��U�t�v~S*��R�L(�y�}���	�m��RP=	PrH��i�׻�;�N�cP�wüA��+�L�)�{rH��i�׻3�����Q�wüA���ȍ�)0f�f�G$�Nt�6��HHD�u�\�Bak�V�|M�̵^�7��߅)�xD����e�> �8*)" ��_Cvi�X;p`�{Ē���\r���㯄j3#��.p�|�B"��D���pa�����Ⱥ=��20{�(m�/i
�\ }Q'(�!��=k�Rm������ g�Q��Ȝxڣ9�$���L�tD:��@�WH�D�n���N�<�\��=�{��M�<"vdԬ��+�Ѩ�f?�R�:��er?G��� ��=����2O�Q�#�ͫa���I˒��M�H�ڒ�9a�	�+4D@��O������݄���'٥��gVا�˓#����!��#��q9+t�}Ż�&ǥ��a���F�LFC7�5$�)�vx/�k
�SR�w�o�FAMs�K-�sǾ�����D�%îqs�~gr�%qV��˚�b����N,���5B�Cy�lj��
�j����H�A���������KX��ik��dc�@z�ׅ�ؘ�X��WG ��@�\����Ԍ��Ǐ�c���w�I�7<�	+�	�u@���kJ���af�iβ�=&��]
���b���M��#l/����1��X��WG ���ָkd�vu+�vW�
�n��뾦��"L?����x�X�ڹ:?�#�6�f���L���ݾ-/�uu��ڿ׏�����M��ܐ�}�q���C�(n5j�?�T���%��X����!Qr�g?	��o3t��F������ӮvZ_��b����������k]���;���h_z�z޷S�xo ���uS ����ߜT��һ���٢�+�����_�˞>��GQ��&Y��V�ٕ����Ԍ��Ǐ�c���w�I�7;�y��a�	�+4D@S���O��zB��݋�^aw��Xá%��v���\�G�����dc�@z�ׅ�ؘ�X��WG ���g24�H���}{5��['D�C�k�a�	�+4D@��/�ciJ�� *�P���Ga��T�rs�(�̴Y�{'%s�6F���y�q� ���+�6e���mn
V~$�i��"u�rB�0j�䴑f��6�k�*x$6�>��?&��n
V~$�#�(pᰓgZP=�����p�>�q�M�4�(��o/���֦N�\��q�l@���w[�>ta�A?:ϭW�Y��RUc�q:�����{~�o{��:�f0u�&�i"&_m��n��0=P�������h�T�JDn ��a�'���*T۳�͕��Ĕ�.p�1��zB��݋�^aw��Xá%��v��c�}���Fo|k�LbT۳�͕��7���.L��h�T�W��S���c�Z�~rw�&�z<aSm�6��`4�04�jf�5ߧE4��Fi��|�3;c�<�o{��:��_%Dό��סزN	��!Y��<YP�pg�h�j��SdZ4�!��Tӧ~kU�#�����1��X��WG ���q�;�Ӄ��g0?��7D�EI��o�D��%��v��7���.L��h�T�JDn ��aP�d�����$�\%e��\9�oA�d��JXl'�&�P�2�PUг�|<Ѩ�f?�R���%\��o.��p*����H��efm�0z�cUL���ޤ�Y5x���:����S�>�3�� �fX�#A�H��~?R����I�
�2�=�@)��۞h�G�jryX2�uso��%����,����«?�z�3$Ȋ���yu�R*E���&�Ut�\�\�,h���y5�����$Hm�wS�$�X��wlT�o��ڍ�a-6�Da�q�;�Ӄ��g0?��7D�EI��o�D��%��v��k�J`�\A#�ͫa���n�e�[7
$B�>���I����~u�o{��:���m4��0�g�F}kQ1�8BW�R7��� tN�y5�����$Hm�wS�$���	�QTXP�e�gA#�B��-M�O��~��c*o��ܔq_�pk��=��hX��9�{���J�s���x�ԉ�>W�{OEׁ��q�2��Kk:)���2��D+���4Y U�����p�zB��݋����f�� !# D���\�G����s"�k
�5��)�rbJ6�~��JUJ�s��\�x���g��̙(�j���%�z�J���o{��:�N�#�@j��{�`��ҜcZ�����c�Z�~�c*o��ܔq_�pk����2%g����<-��ic)�̩��x�ԉ�>�e��@���=�����Lj1���7GX�=1�����
�^��j"-M�O��~��c*o��ܔq_�pk��=��hX��9�{���J�sׯ�ɛ�?өW�{OEׁ��q�2��Kk:)���2��D+���4Y�q9+t�}8BW�R7��� tN�y5�����$Hm�wS�$A�~����9���&�޽Ut�\�W�{OEׁ��z\�Q��TXP�e�g�6�<+s�q9+t�}����d�n5j�?�T�LW�_����V�&ݡ^����;q����}7�������\�2���.Z��'���:��KY�[b%Ɨ�W�{OEׁ��z\�Q��TXP�e�g�6�<+s�q9+t�}����d�n5j�?�T�LW�_����V�&ݡ^����;qf;[���rw�&�z<a�4�ڈt׏�����MB�R���>_Ѩ�f?�R�Kr���щ���ӮvZ�k�b𓣊���%< �A
��z(�����N��۞h�G���=�,Н��j���J�������ۧN�g�c�`�zR���b�S�w҄���m�c����p�^1N�����T��E���q_�pk��=��hX��9�{�� �ދ��kn5j�?�T�^'��s_ㆂ`Z"�AJ���U��Ĕ�.p�1��zB��݋���>?���{��G�����
�]W0�e ��Hp9���o{��:���m4��0���f��J�a$�Y ��\bʏq�2��Kk:)���2��p�!���׏�����MJ�1���۪	�}a�]�w%�oφ��<�6�w�i�����������)9�1v�1W2��,t�ZR�F�"5�Ϡ��)�\ߖ����-���ZA}�/6�o8:4����=/�F�����ٕ�������=/�/�� �gj7�cL���	Ǹ�y85��*�Vy92_k-f��%�n
V~${���up>'Ίѥ֤�g�-�Lo�{ 4a��|�&۪	�}a�]�w%�oφ��<�6��B�Ә���!�`�(i33��0��7)�0�1�!�`�(i3M �̦�P�c��f�.E!�`�(i3!�`�(i3M�!6h��sȸ�"rR!�`�(i3���S�K���Fz�!�`�(i3C��F����]�U��!�`�(i3	Xv��#E�l*�����l*�����l*�����l*�����l*��������~q,�	iV\bւ���-r�_?!�`�(i3!�`�(i3�Y1f��������!�`�(i3�6Y^6ь���ݘ
4D!�`�(i3*M׷��!l*�����l*�����l*�����l*�����l*�����5$�h�Psȸ�"rR!�`�(i3�ng�[�^�6Y^6ь�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��5䳽!�`�(i3_j��u��[2�����Vc�/!��v�22�����Vc2�����Vc2�����Vc}l���fsȸ�"rR!�`�(i3�'e��Ď��`�h���N!�`�(i3x���'RFt���g�!�`�(i3��5䳽!�`�(i3_j��u��[2�����Vc�/!��v�22�����Vc2�����Vc2�����Vc}l���fsȸ�"rR!�`�(i3ɦCNM��FY��/׷�n��`
HF x>H�|�,*
���i!�`�(i3��5䳽!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�&E��sȸ�"rR!�`�(i3!�`�(i37� ǚ�y2�����Vc\�29m8l2�����Vc2�����Vc�inca߫r!�`�(i3!�`�(i3!�`�(i3�x�?J,���O*���=�����Lj%"d��&�sȸ�"rR!�`�(i3!�`�(i3�6Y^6ь�I��&� ����ֶ�!�`�(i3!�`�(i3��5䳽!�`�(i3!�`�(i3!�`�(i3��2}O�����:�2�����Vc2�����Vc}l���fsȸ�"rR!�`�(i3!�`�(i33��0��x���:n�q m�e���b\�#�\�'�ڦ���X��i)��]��ⅴo=�I�r�I�τ4��3 h��7D�EIdQ�;{�r6]����ez�:Y����"
�����]�DP1Tb ����IX0F�M��LV�!��o�½X5 N��r*<��=���jl�iYX��R*E���&�Ut�\�P�<��^NE�g�������(ӈ��Z��&61����g�Z��3��a���Cوj�~Ut�\�f�hj�"��Ck�8'��d+������1��X��WG ��Ѩ�f?�R��f�;�>)�-��a�A�([��}qn
V~$Ѩ�f?�R��o{��:�N�#�@j��{�`��Ҝ�@`��@��R*E���&�Ut�\�Ѩ�f?�R�x���'RFtI��&� }iIB?�j�&D���Z鎬�������(����ЊҼ�<��L=X�� �-M�O��~�����m��^��dx=]�Ϲ���6�|�MX�	��*�kv٥P5���rs�i�Ǘ$� ��������-Y(��%W>F��)�_�� Y!܈��u@f�u\���:��΄x�g��	��S8��<��Qʵ����tBp�l���P���ү�+ҋh�Qf�
^����݄�����;R���AL%�jvo�HT蔊�cٰ��]�Ϲ���6�|�MXj��R�6Pih�Qf��5ߧE4���q�)]Q�x��r_��m�i��"u���Ȇb�L��B bb���H��efm�0z�cUL���ޤ�Y5x���:����S�>��a-6�Da���˿1ϲvv��I��DЎ(��rs�(�̴Y�{'%s�6F���y�q� ���+�d'{���o%�RL������ʵ�����9�W�"7�cL���	Ǹ�y85�΍y� I�Mkm�m#�m�e5ngY�-M�O��~ӶC$�-��xM��R,�g�zSB�������h��}�mT~1�����(��(����ʵ���ه� �4�<rw�&�z<a��r���x(�i��/RvE7�MWO�6�c��$1ݮ�I�C��,�jK�3��u�!x�R���- ����%7e6����k�'�d0�(_� gg-	�\�G���:��er?G��g��ǻ�Ji��ċ�!-M�O��~ӿzR���b	;��Ǧ�<z!N]����Y�1Uj�|ᓆ�~_Nv���å;���.[r�gc�JV����l P�7��Hn#������Uh1�z�X
3kZ��5ߧE4��p�-a�D͢fU�9�׏�����MFi��|ր���5V��	��yx�_uE:+4����_pQϧp��k�����z~U�6B�Ba��;>�G]�K�Sb6�A�e�r���b8#۪��������`Z"�Au,���Ex���O����_��s�֙P��gg�@��uF�J� D�ԗ�CW	�h0^U ��ש�F�3h�E-�;�]r���.~i����[��%aWp��.�替��+���<j��ʞ[��;+�sb�]��A?�X!�2YLވ�]� 0��CdJMaM�Bt�0�:D�?��l�����h�x�(��d!�!A��f����$7EUf���@\I�r��r%��ό�;�LȫԷ�/ᮽ�5�"t�20{�(m��M��X	��!Y��<YP�pg�hN`K�7�I�b�&�q�2pn��gn|�P� &G�N�g�c�`�ɺm7�{�݄���K7͍��|��W&":t���3�l��d��JXl'�&�P�2�PUг�|<�D�$0�y�R�QY`�CgD�|A�$����@/��r �a�<d���u�q0O�*2t�ch���5�����Qa�	�+4D@vE7�MWxM��R,�g�zSB������ɲF����z�X
3kZ�
^���cv	�-�?x���sM�а5�c�ؒ,�X�nrm؊(��L~��h��3K�<�
]3b�J�X�H�u�q0O�*M��3�}�v�5�����Qa�	�+4D@i�a�sir�]��<�A�FRsyѳ�)�5�F�Y��(�-����$[���	x=:����fd�P�<��^N,���}a벩��Y�^~>��mJ�1���K���L���4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY�c����gp��T3Z��	�J�-D��`ʏgG�H���b��@��` �6!7�_%Dό��סزN� �w���zF������?M>��^J��3��a���Cوj�~�4v!4���u�q0O�*M��3�}�v�5�����Qa�	�+4D@[�^�2�f���jv�':�j��� nΗ��FU�D���9�@�r#�9l$U̑�1G`3n��:��P��Y�K�4���jv�'ݟ=�NM���\n0�8�׏�����Mx(�i��/R�������a�U�ے
\���1�k���^�_��r�I��oI�u��qAxDp��T�/i�M������t^���\�}�]��Ko��M��X	��!Y��<YP�pg�hN`K�7�I�b�&�q�2pn��gn|�P� &G�N�g�c�`N5L�`!|�l<�K�旼��7X��^w�̀�l"�sW��/dN�<@Iv��nt=:�z�X
3kZ�(w"<��J�F�Hj��b_X�XV�b�z'hۉ)��R��삍(�V�ܼ������A �k+Q�h'�Ȝxڣ9�$����3�� �fWT
Y��%r9���TLB������([��}qn
V~$8Ơ4�ܩ"۞h�G�2B�_p\_R*E���&�Ut�\���x^+�����.� U�O��5��g�g�D2�+�ܰB৙��7�0)�kEu��-��e�=G<7�#�z���f�DWogyV���ҡ����a�#�ͫa���n�e�[7^�,1�NgWaU �I�%�z�J���h:h_Q\��i,��fx�W��L�7�+fqQ�y*ط��wƑϥ�g7U\a���5Cc�}���Fo|k�Lb�\�G���Wxxܤ�]
���b�v���V�i�;�H���o�4�= w
��ݔ��������@/��r ��%�z�J��A`g.d�q_�pk����2%gY0��xeð��Th�Qf��,2�C�����d���Ą�Ĺ�,7�cL���	Ǹ�y85��֟��D�D���P�ħN�g�c�` e8�~��Q�%q�E�����"��C��D2�+�ܦ��)f�V(��Q��\�ͻ�.}y��@�piM�k}���u���5������ e8�~���,2�C���l�yi��L.bC����������}���u�}S��Hō�a-6�Da�l"��Y��WwOkd��l�\a���5C e8�~��(w"<��J������!��&�i
Y�M�<*LF�#P�j2E�?J�1���#P�j2E�?T۳�͕��4ޓ���@l��l��n��=���#P�j2E�?W�]:vx��3AE�p|�/�GT�)��3Qk�	��5��g�g��)�-9�4r��g2�~��R�MI���X�=1�����
�^��j"�*#�IQ܋����� 7�+fqQ�y*ط��w��c�{rS�b�8Z���%\��o���h�Me!d��q杳/��-0��3t���=�4�04�jfu���%�[�2Tƭ��q�j(�+�}��ɣ8��9�.�`���c��u��-��e�=G<7�#�z���f�DWogyV����T۳�͕��9�d�L�� *�P�RO�?@Pf)�+�9-�i"'���Xw�j�7��FZ����^��h���LX��WG ��4ޓ���@�#m2�~�PM �%�s�~����gyԡ�U�y���\��2�ĭ#�?UM�#P�j2E�?x(�i��/Rh�Qf�(w"<��J������!��&�i
Y�M�<*LF�#P�j2E�?�5ߧE4��c�}���Fo|k�Lbx(�i��/RŻ�&ǥ��a���F߸��S�Ȍ��"+VqS?�d���&����I�����^�_���=-�!�^G�*$\���/�\U:�aw��2V�RGS��=[��uܖ��m�el[������O����_��s�֙>�5�(2�q�is��g?	��o�dEr�+��#ȕ�B�������Ѩ�f?�R�g��j�([��}qn
V~$�UӇ��ɋ� ��X�D
CvK}D�؈a������h:h_Q\�=<�6>e��0�U+�qbp@�p�-a�D͢�����.�����T��6\�4�@���(�?<n
V~$_�)!c���~?R����I�
�2��.���-M�O��~��D�$0��5Ɇܾ�]��	He$(�2�ft+�f�;�>)�;��e~]1bt�Z��P��3�Q#� :a�	�+4D@i�a�sir�tFy��j/�GT�)�[�=�({���*Ȣ?u����E	E��D�$0����{?tQ���WYG:�rs�(�̴Y�{'%s�6F���y�q� ���+�6e���mn
V~$�l"������3Y����Q����ۉy�T�����j�ew�]����z�,�X2��3t���=�4�04�jfrw�&�z<a�4�ڈt׏�����MJ�1���۪	�}a4����@[�_zβr��S~��d8i-9���a�d�Ĕ���e��cx��K�XXz޷S�xo ���uS�yQ��b��������Rܗ_.����������l��5�9�e0���0��/�1��P����^_曕�!y�����qtn�4�rxE�N %c�G˜�}b�J~�ʒ�B��u����&����~���j�f�o~��������,��j���a��d��t^�����P�5��t,�'��.	[���,d�iл�.��L�u���X MY��w�ܹ�YL`�Þ@_+h�J�}���(w"<��J��Ȇb�L���v���Y�d��&n�O��0���Ȇb�L5$Li�E�4{�}j� ���ʵ����Ƹ.��v�X40��7e0���0�]T�����7��<�DK�/�1��P����^_曮�S��%[����;���~��aU���.�h��[C��ԅϪ0^�j��WV�#aطR
�^0oߙ�(ml���d�����7��|�K������_6j�"HsضZ�i\���ޒ�#] 
���8��pP�ʭ��2F���rcJ]�0�6��b�gi��#g�k��΃xI��o���%\��o�݄���r�gc�JV����v�}�h�]�V��t_-Z���Uh1�|�+��?�d���&����G�٘�&�T����0��g���>�HGt���/i
�\ �D������V@BɇF�����k�O�۲��[V��M*�&T��L��o���wu6�M`B�Ӑ�>�b��O�=7�}|��	f��{#�~��:����嫋�T�%][��"��0�ʂ�j�Ï��	�Li4"�	��z��R��/i�D�]
���b9�s}�T�s=�du�([��}qn
V~$��D�a��^���f;[����w�򪥃.(=����5۞h�G�jryX2�uso��%����,����«?�z�3$Ȋ���yu�R*E���&�Ut�\��&�(5�;2:��er?G��g��ǻ�Jt�Z��P��3�Q#� :a�	�+4D@�K:+>�Y"�g�YZ6��HHD�u"�T�B�Z�R*E���&�Ut�\����˿1����{?tQ���3E��٥P5���rs�i�׺�� �������-/J�����Ut�\�Z$R�Z�]d��l����v�}������Ja�vݝh�c�A�L'B��o彍/Üy�a
��ү�+ҋh�Qf��_.�������0=P�������h�T�JDn ��a�'���*B�R���>_r�^�#v��.ȅ��J �ҋ�;#P�j2E�?�5ߧE4��c�}���Fo|k�Lb�e��@�;�H���o�����jw��1��X��WG ��Ѩ�f?�R�Kr���щ���ӮvZV�Wg�vy�R�QY�v��|���@F��ɥڦR*E���&�Ut�\��i��"u���Ȇb�L�($Z�u��΄x�g��	��S8�M�����vg����PTse��ͳ[�%�z�J���!���睋\��@�E�B�f��.�zB��݋����f�� !# D���"L?���C��׍�߃��:����嫋�T���Hp9��x(�i��/R�P�HS|�4�04�jfJ�1����ݾ-/�uu��ڿCt�w#��@�������a�U�ے
��7�j�-!�7���X���סزN� �w���z����T �o��Ow;t4��(Ic��+h}J�z޷S�xo ���uS�yQ��b���:������p�Ԟn�ʚ��^�8n�G�Z�Y�'�Ԅ�F{����i��&�'J��^�Gߔ�M�t�5����3�����Qbݙ�-M�O��~ӎ;�z���ΥT�t5IйP2��O���ˎ����(�?<n
V~$qSm�G۞h�G��0�=��l��j=/x9��g��ǻ�J�H�ڒ�9a�	�+4D@��/�ciJ�Kr���щ���ӮvZ��S)�3=7�}|��	��a-6�Da�zt��[��T�卩 ��������w�򪥃WT
Y��%r_�1�J��]LB������([��}qn
V~$T۳�͕���\�.�ϗRأ؛��3Y��P4�a�?O�0|��ˊWKkH��g����Xu������6���Lv"��D�$0����{?tQ���3E��٥P5���rs�i�Ǘ$� ��������-/J�����Ut�\��i��"u�rB�0j�䴑f��6�k�*x$6�Ú��\�iUt�\��4�!���];�σ�������ng��	T�B�R���>_J��}0�^�s��R�����jv�'x�W��L�rw�&�z<a��r���֒.�N�l����旔+�ez��2���թ�~X�D�����+�=�b �\��)JT��w�򪥃]��9��6���ʵ�����9�W�"7�cL���	Ǹ�y85�΍y� I�Mkm�m#�m��h���LX��WG ���"L?���J��}0�^Jq�l_N�4F�sltPM �%�s�~����gyԡ�U�y�z�X
3kZ��5ߧE4��p�-a�D͢fU�9�׏�����Mx(�i��/R�������a�U�ے
(㷾����[ �����
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.�	g�yߑP�~�I��~+�.�Ҙ磋��w�����H���D���0m$u��+�����oPJ�F���s�V�����Y����딼�\�vūx`��:�֡�\�<7�X�e����yM��$��XP��ȭ����m�cc�PƐt
����������\�v��Q���K�1�����C�[���Q�#<4^��o��C!T*�q���U��3s]o?�E����F�ҋX����@�ڗe'�f�;�>)��U֔�>V	�]�!��	Ǹ�y85�R�m�.wa�Iz#1�<Td��"X��[���1��"8U#��L��H&���'ʤiΉM��s�>P�2-i_���F��
S�>��Z)�� ��P�$ke���FW+w�7�jU-j�`Z鎬�������(������ Z�U��c-a(􆿳��WakemDK7͍��|��W&":pzl��a�$I��h\7s�9���o��S8�[��>�%MM
��,=(���4ܹ���fNd��"�A�S[W���>V+��k���0�:=��C�Q\%?D{�q&�wȽѫ�	|�yv<�1���\�۟�-?�d���&����{ԕ�/�����jt���@
�ѻ��`���+=����7�>D�c�lQ��� ����7끍J�[T�)���� �&��׃�`�n��U�z��pU6�M�S��2�{��΂�W,x��k8�5�>�yKYQs��[�|�F��ˮ�pd�Zз���\��6�R�X�?�I��H���Ku U�zjb01
�;��S��y9Ez��}��H֞��� �z��w�����4L"炡t�8j�t�Y�Ij���0E���FZ���;D8���:��M�S�ᳰ��X�z���t���Xo޲G�����$7x�c >��}f]���]�w9"x�g�Hz���MN����!I/�������A��1��+�W�Ń�I��-NdRg�/�mC ۸���9��;9k#:̧�	��U;.��=IN�������ػ(z��Rr�kB}'<� �w���zF������ݚ�Н��df�L�_dj�Ï��	�Li4"�	�Οe^��\'�s�@#Fd8�^S���$I��h\ӗ��= �*!�`�(i3!�`�(i3!�`�(i3t�Z��P���]�K��l�u�;�A$������l�u�;�A��h�S�~W\'�s�@#F!�`�(i3!�`�(i3�7-�^x9%�fu�A]���� *�Q�駫�]���� *�o�v�ԇd�c�(��t�Z��P����磱(f�Ah��p)	Z7��Y�X؝�h�rr�����Nuv��b�0�����Oam�.�H��`�M�ͦ�J {�ú�8�$�N\��
�Mn�Xl`�D!�`�(i3!�`�(i3�it� B��@֗�0
�O���G9ziJ6��7,ʽH��L�}�oW<���"��Тϫ��8��/v.V��T��#�-�p�������?�r�J�2E-�Rxp���[0��]8��"��Cl�3tu]�MP��br6���:��j��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�k�X��0М;�N�cPkax��.��m-NJ�*�6-��9���v�)�BҺ�)�|�$N�?��N��0��Y�b�0$����!�`�(i3!�`�(i3�%_Z�ք{q��#�i+����Ó�#��d~�/�3> հ�`�H<�b���ˢYۋ!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����k��J�Z���>H��L�}�Lqo���"��Тϫ��8��/��X�˾�c�#�-�p�#��d~�/?�r�J��4�= w
��D+���4Y!�`�(i3�����L�	u]�MP��br6��ۻ 288����Q�U��Dٺ&�Z�Ӻ�ew�T'��8��	͂'�)������Lqo��!�`�(i3!�`�(i3!�`�(i3!�`�(i3rz��G�;����A=&�������*�yȩ�,�=�'����M�m-NJ�*�d+st�I6�v�)�BҺ�)�|�$ h�-j�(!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{�[��E�p�`V�xs��4�= w
��3> հ�`�H<�b�uu��N�B!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�`�>'r�:�;�ࢄH��L�})��yG��"��Тϫ��8��/�v���V�i�#�-�p��4�= w
��D+���4Y!�`�(i3!�`�(i3!�`�(i3�����L�	�U��x]�i�A�Q�8�:��j��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�k�X��0�k��=��kax��.��m-NJ�*����6G4ޓD+���4Y!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{q��#�i+����Ó�p�������3> հ�`�H<�b�N�)��l!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����k��J�Z���>H��L�}����Z�"��Тϫ��8��/����BSb�#�-�p�p������?�r�J��>Uv���ߓD+���4Y!�`�(i3�����L�	u]�MP��br6��ۻ 288���ߥp�dyeݺ&�Z�Ӻ�k�jZ"��8��	͂'�)���������Z�!�`�(i3!�`�(i3!�`�(i3!�`�(i3rz��G�;����A=&�������8(<���=�'����M�m-NJ�*�%���d��G�v�)�BҺ�)�|�$��Wi����!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%_Z�ք{�[��E�p�`V�xs��>Uv�����3> հ�`�H<�b��<��K��w!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�`�>'r�:�;�ࢄH��L�}�gÁ�r�Ѩ"��Тϫ��8��/�7e���ss�#�-�p��>Uv���ߓD+���4Y!�`�(i3!�`�(i3!�`�(i3�����L�	�U��x]�i�A�Q�8�x(�i��/R�������a�U�ے
X�q�	��ؿ��=�M��0�d(_\�^?'qKy���\N}zp�jN�!O�1�xI!��6$V����W�������9jx-Հ�ue'��ǩ��or��	P{�R�$�V֟����J�FZv�,�+�]
���b ^�x~�(vi�t�c,�q����Uh1ݰ�:l���K��<�Iz#1�<Td��"X��[˽�����3Ah	)ޟ��E.t�