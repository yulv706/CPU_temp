��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�Jз&�6��`�,�2����yׁ @'�إ��(�q�<������0T-~�	�Y\�������/�'o��Ӻ��,Q�Q�?uG�Qy����JN�YQ���b`.�]2'%Sǘ+�����I�'�z��9���
cC��O�-��G�s���R����#1X�.ՅT��+Ϩ1Q�2�:C�.0q1��B�ce�jͻ��}�����9�Kو��. z��ڠ�1p�W��b࢞�i�Ot���k`��$r�^�A%�7��� ��R�āy����yoZ�P/b^��GAjc*!�� �]K�lh��.��:H�T�fޮ��Ĉ;��~h��h�W��>�:��)�򹉓��#�)��#�)�� A�}Z�n��-�4�E͉�-�DfWn~��7��+�gE��e��d*��N���9׬��Lw�E*��+.3����sv�RS�6�1M���yK����ॶE*��+.�}���n9��W�Mށtd؈��k�;4���Fz�	�$C�jQT	�$C�jQT��x���t���R=l�#�	�����g�Έ坩� <�44��v��,X���.�bI	\����	d�ዊ}��~:�u���n9��W>X[V��k"Y��^4~B+�9�'���Fz���Fj���Fj���x���ti�8P�-�׭{6V_��J&���1�c�ؒ,�X���2���O�hf>Ŋ�g��@���"�Q�8t�s�0���8��t�\����1�x���0��%C��0̉YaA�=̮Bq���'�y䜠�:�A�}_�r�t#�+��O��oy��09�nXm:m�t
�W_���1�o��Sl�xdG�!�5��� ��YY_���6�z�
^��1���K���π�>���cl8)��� ��J��b2�K\��$����\O%���F{�? ��:��c�b����f��Y�5�7cWr��
�1�ِ�E㟪g�7�������0A�OT<��y���@��v�m�qs,�Y[Ն�l��"F6 崭��oes���$q��mKx"E&��� �$Y��C��s7Ҹ���/JF[B����,q�.3��h�V�*�U<������P�S�bN��4( �.x�����fg��ͥ������QH�<�h�d���@빮��1o���W+N��<�DU]sȸ�"rR!�`�(i3VR��|B���D���
�չ	L~�BA�kN��&94$2�¤}l����Fvf����P��~w����+���m@�p�Y:
�B'���a(G����h+=o���&>�S�䡢��k͝�ul���C�A:���i�����Fz�!�`�(i3��^�j��VR��|B���D���
�չ	L~�BA�kN��&94$2�¤}l����Fv+�-EP,]�!�`�(i3������=O�Z�:���ro�؛�36�ZpMu�IRIn����\'tI�D��ܛ	g�p}XR6��^U���Y!�W�Vc�sNL�u�
��Xx����G�$�-7좎E&(p�
����d�k�ViR��W�ik2)�
}wʭU&H�1��8�h7H�u�ÍeZ8��
;��d��q�G�a�P;m̳�UlgRQ�t|Y�f�sJ�F���s�V�����<o�nïi�JHn��z��r9�3,�qo�,ܛ�	��|��	(���zL͊�q���b�Kzb�d&(C�#�7#^�Vn�^ֻ����XP�����-����[�f;q�sɈf�=K����X���`>;�`w��^e@��V��M�P�zL͊�q��o���.N�wJ�G�����t �JHn��z�w٩L7���i�^e	�F�K����'�Z������be�o
85�C`+�9���m@�p����
��s6��\�v��wc�}�![W ��"vY0Jߺ�'n�^0o��]�mj:�ǆ�0��n-=1�BF�k͝���<���r�����z5Ā�����^�j��C �H?�o�ݷ�����.j�,�3*������|���kJ�|��].��'���Xw����l���(���e���!n}y��Y�{'%s��.|Z�����@	Q^�V]��}R�wX��*��p��U�d�K��@�!n}y��Y�{'%s43u�R��}/A;T�c���Y#?M��^e@��V�m�C��x�T�\ ��fȂ?�x0�C�Z���8k>6s����]�!��$��lW�d&��b8��)R�v�w\�L~΄gO�3f��*����f���,�LoG�ٳ��?T�]D�9�ϑ��[��;e7�)norǟD�uiL${?�����>��yܛ�	��|��	(���zL͊�q���19TH���'�3�$ �#^�Vn�^ֻ����XP��Ȼ4�t=�j�.�/'�����W;5B5Y+� �i7�sp>�O����!;�Y"f��g�o&�Y��>�_���ˍW�}�ke�Ts
��q{�f��a�/������#��=ό������?*	�ML�벗0�HC�a*�u�&� LK�a�]G��wi�bZ��b�Bv�~������]�!��%��rSe�u�heJ��Dv�~������]�!��ߌ�>!�0ӆu�۲.��!n}y���q���U��@���Ϧ��Ig`i�ҋX����@�ڗe'�D��/���_3#ڸZ鎬����R;j?�鴜�֞W��{l�f|�ό���.�c�{dϨ��B�>�9�6�vg;Je'���Xw>\��p}�	��D܂�A݁ؠː� ^��y�C�9a<�YVKsz�D�W��Bc�i}3�J��؈��k�;4��K�Q8@"��_o�'�Sx�lޞ��rs�i�jf� l�ǉ��F1x,0=]^	�&������$Y��C��|4�ȟ�|Q�P���2��d�٣��c�A�L'��!�a�&H�[&-n�g��U-�e5��e6²W����_]g��
F�UTz�`�J�'���Xw�j�7����ӳ�Y�
X��������`y���pzl��a���#�NN�y�����Ӑﻋ-�����S8�/ #O�)��BT�^��a(􆿳���L��F[q磫��<�:�π&KXҷ�YdS�=��6��+ͻ#q�H!l�5w"^	����3�K���蜍6���Mf���9��Y�{'%s��.|Z�����@	Q^�V]��}R�wX����K�Q�LP.���.�D�m �Oh��M�aQ�q���U�pzl��a�&W4�b�A�w���, n}]�}��V'���Xwa'�<� \��5"�7t�J�4Is*�I94�0.��=Y��_�0z�cUL�%*��"����A|��`y����s��d�\��MN����!I/�������A��X�@�5��6�l��s�����[� y�~��ż3���F����T�O�H'�J�����=<�HI����>�W�_=��0���̏�u�=Cm�v4��61��7a	�����Y�
ɸ�oƴd��t�'��9ܛ�	���V[�+
�l掝�K\m��U}�	|^�׽R�s�DH}�_z�9�E�\����8�i�`!31u{w�S� H"�nT��z��uWU4y5=>F/ġ"���Չ-d��r�b+ӄ�bİ��i+��*�I�GIN�|L9{�U���-~M�n����x5=��{t_�sVh�a�ohWt�_a�1�܄:h	}4���!�fJ��l߮�pd�Zз���?̕U�/j�g4A���{0Yafk��r.y����nL���~C�V�T��a׈Eg#f�z�q���<�{�!���"4��:@��o���KEd��]^X0��
x-	���'�$HgL��)������e��Q�Q&I`��=J'����r
���I}}3M�C,����|#^�Vn��l�M�c���=^��>D�c�lQ�����+�7끍J�[T�)��o�B��^�֌���<�a)�m�d�so�}a�C�ub;�;���dMb3���y�z�ۼ��uWU4y5=>F/ġ"���Չ-d��r�b+ӄ�bİ��i+��*�I�GIN�|L9݈u@	���M�n����x5=��{t_�sVh�a�|�&�#�E�d���������|��=;��|B����?�IX[��O2 7�,�)�C�BS��g\��ı�ZnZ���qq�c�@,��ڬ�A ������ĎɌ�[9�-�Ҧ�{b�J��@��$L��%��Z��b,�0g���>a��v�<�RohWt�_a�fC��0��:Y����i%��ό�;�LȫԷ�/��Ϥk�;��|B}ø��y�w8#�RC�G�G~��6 ���F��G�z�e�3�ԳN���#t����n���n�".�������ܫ�o�k>8ih���A=���R�O�����m@�p�����Ш;��|B�[�%��PCd}��c��D�m �Oh����V_V��!Z��|<;��|B�����m���6���s��y9;A{A�k���>�*7�=�6�Uw�ѥ�+Ȑ゚�H3�rwJ�G�����A��9W_��s�֙��h%��i��؏��=O���[�_7��ҩ���*���6j�"HsD�A���T�o�k>8ih���A=^��ܑ0!yN8���U���-�?,��/T}��]�?�y)�x�d��cɁ#g�k��"����J�=O���[�q� c���xsq��?�d���&�&aD�4�LP.���.�<\�9;L��૵�`MoqF}.	�jo���wJ�G�����A��9W_��s�֙f�P_�<�ey;���W�b�aY��m[�c�Z�~����,�ǰ�.��յA��Ye	y;���W�b�3����|7�Q��wR*�e��Y�!��5�q�^��𔜆�x���� ���Qo��#g?	��o�ܶ�p�2���\T��y;���W�bx�E"�i� N��r*A_��	A4��4��Ǳ߁��BT�^���8�B���A��bu�x���S.ш0����be�o
��sd$2�,��$f!ٻ"�%2߸��H�D��=���#�NNҖ׳M��_���"�׼L:�%��9�]�3����s�]�<ܥ��QE�4�4/�c5wU2K� �M�����<.A����8@"���ⵛ����X^W�E�eN�cb�e��|4�ȟ�|��m׸c��V��$���Y#�5[u��Ƴ��^e@��Vz�+ʣP�S�8G}/Իj��&$�^��V ��������b���`��f �̵P�B-�\&A(`#����c�Z�ٹ!5�j�BEޥ�8{��o@)�A�|4�ȟ�|ֶ�T=��v��z�(Ԭ�����`^�	�S�_���k�:�j����(�V�ܼ�ʽ��φ��<�6���k�J��W�w��fD������Q!5���`�(���}��vt��@�mǀ�A�,#6:������`V��ˀ��u��6+`O?�Sկ�M�[L(,�$W�Έ�:x�����诶�|��:��Z�j�t�R��A��E�5�?].�`�ny�;�>�=H�����0�]'3�d����l�F�<����I�+ ���������ĉF ���^3O��IZ0�s����S*;p͊<^�D�F�����Z͝�O�~��3���~�8���4$6EQiĂ��*����ѿ��Kצ[��EEp-�.�^��K�(����q���d��^�d�}|c�q{�:/���)�������aW��2|�������XkN�U�@Y����!|~��s�;�9U���JSo?�d���&�G�`͈K�Ӧ{Ԭ��RA�q�m�,&H�[&-nD�P�E6�k��q��־��)�!�B`�M̛��o��o�iCorǟD�ui9�f?Y�O�D�c��QԽ�>��yܛ�	�������,����|#^�Vn����a�:�n���������W5�\tCՙ��BC?T�,����_\sQQF�;�?2^�9<o�nïi��n�5�F�^hq��:�����S�|�)LE�?�y)��0�sfPEwJ�G����������?�_��د��� r�����
L+���N��7�ͭ�s������Y=��~<6����K��J<W�f�ӊ[�k�T�"2o�I���6�*��!���α�%�����h�f��Ҩ�_E��ڒdk��������h4c�LU46�0�� .E�����ͮz�w�	 ����h4c�LU46��>��Qp�U����x��ʢ��ch���X �8@"��U���F����ۧc��U+���(�uÓ�h;�.��X��!{��%31 ��e��蜍6���h���R��*1�#�;�N�ߋ��[�Ee�&��c�����|�\;͖����,�ǰH7"LTft���U�2����q���sM,�%�H�n��шI�֟����!|~��s�;�9R5Y�4�;��|BDt�e�v~ף&��W�4��Ǳ߁��BT�^���8�B���ow_;O
�xkx U�_@�Z&)������%7f�=�٧�\�T����!N�~<6���xՉ�T�Ұ>D�c�lQ�2�G�Ml�y �谝��X�e�6<�AT];�'�3�$ �#^�Vn�����'MRmHX���y�XZ@po8�.�V���c�PƐt
׫�J��!��l��[�?2^�9,����_���3e%��P�S�bN��P])Ƶq9�+�ty��@qW8�e�Ts
��y��T#¢�7@�@-0|���1��P��gΐֈ&����|���kJ��K�}i��$�*$`��'Ƶ�s�(���e��Q�'`�����-Wi��'�㉨��ӆu�۲.ȑ��O�v�E�>��w�VI�a	�㉨�����D������O�v������%��{uMѧ/~�9�`u7M�j��LU46`��f �p�U������5��\��h���X �8@"�ѯ�Pv9��A���:kug��?`-ʂQ��RU떐q磫��<p����,c��%g�j�ym1�H��ۗp���x@[�_zβr�v������]������pD���㖄~����ptn�U�_%,�}.ς�n���㔡�ʁ�;C��UѦ��	}�J���x+l�utO���!�nφf��B�o(�bkֈZ��h:ҹ���7�K��#\����s�;�9U���JSo?�d���&�D�;E��D?�nϨ�_S$?���S�������o�J��p�a*]R���ZHOh#�×VW���(��RʹZ����Q6D���WX��y�g��U-�ed��
���V&(^�og��?`-ʂ��Me#p1�';��#js䐼�D��4�L^�y���c�Z�~rw�&�z<aSm�6��`�E`���\�ܢ��,a�U�ے
 '����X��m�l:M/��=-���K��Ƕ@[�_zβr�v������95���������Ρ]��_kjY%�4��d����Vu��uz�(�E�������� ݟER�/�蟞w��g�+�Ĳ�6wK�����ø q�M�4�)[9{���E8��]3��&Y��V��E.���?��ʮ@6B��x;�-MMk��*"}�ή\}�~��k/�Rp.$�Z�G�:y�j��kd�5���Q6D��RZ����c�*�&�'�UKA�/6\�/c�z�5T`S.�<�T�V��\��5r$���bAg�
d�mEF��y��Y���q���D�	�$��1�Ч���[��+h W��]���"��J�$��Ϳ�QNJQjO.�r���$�N哄�f��ϙ.����n��݄*���-����o+}���
�L��	V{%�Ӯ C�`�j�T�!_!���U�p�J�R�r��a�B:ҹ���7�K��#\����s�;�9R5Y�4�;��|B* ^���x������������J��B� ��~����rZ���΁�Y� 63��'٥��gV�<��H�HtA�q�m�,&H�[&-nD�P�E6�Εq�8�W)�x�F[*1�#�;���p#���8k��.ͥ�P���_��r/��=-�� �F���%��v��p�-a�D͢fU�9�Ct�w#��@�*�W�Ǹ!2�͞nOY��`^�O�a*]R����]���3Q������iԄgc5E.E@�Zx�L��Kj�9�I��&,Ξ._�0h�5e�|͹*�cW���&Po�tTs�B&���]����t�>N�z�"�~�����Cᣨ*��w5t�}�p���� ��M��7<���Hn
V~$�����lJ�4Is*�I94�0.j~�]����}|�$V���Z�%�΁�Y�ה��+���F@�m`C��8� �����A�ip�-a�D͢fU�9�Ct�w#��@�*�W�Ǹ!2�͞nOY�s���{��9�2�LiԄgc5E.E@�Z3F�c����;�
�8\),I6V��	��yK�)ر}�!rJԱ����A�H1a�k������1��B��m�E�='��9=VU���_��s�����%8���}0x�%ѻ2�ͫ:��e��q�y�r?�R�?ӳ��S+"�{!|��Gu;��4.Mw��\�� {���L�>
�h�7G>���	�+T%2q�,J�l�/,�\�׶k��)�)���a��-B^b`��qm_����~w����+�#���]�D��ׁ�~vZ�c̱���W�k"�f��6��-KW�*�	SE���_�o ��Z�� �s�1c��K�kMbY��X�����f.��2$6�sI�U�z	��v���ܠqJ��i��9Ua��O�H�s��)��7��2�Ζ�7E�'�o~b!��u�n�Ak�������s�]��;*?�|9E ~k�w��!�@MiQb!��u�n�Ak�������s�]��;*?W�J[k�w��!��^饑���b!��u�n�Ak�������s�]��;*?���4 �k�w��!��w��p���
�C~��go�+�Eާc ��$b�[��|��M�[G?�#�
y4�t��+��m6
�DR����X��wd6$�gd��U���A�c!�ܽ��=�z�Y����S��.�����6	oO��z��R(qq�A�3J#:�� <݁&�}���
���*,f$�7Q0- ��Ck�fÜ�2/ͭ���Y���1�/�I�����;�y������,�p���>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z��r9�3+��8����Y�I���^ֻ����XP���Kvq�?C�$k;e�q��m;5B5Y+�T�����N��=��-��5��ٺ�`�� ��3CO+��T�D^HUB�����#�q�£.D,����e!0�K�_3#ڸZ鎬����Ǟ��݈�<�){:�|��].��'���Xw۠̉G����Ig`i�ҋX����@�ڗe'	������|��].��'���Xw��C��T��Ig`i�ҋX����@�ڗe'���'5�7~�|��].��'���Xwě��%� hZ଻|���9�dMbZ鎬����+��4{��8�O�3��ۋQ��T�&���#�{�0;�}� �ԕv��t=�� VU+I��B<�p�@���+q����R�0{�!n}y���q���U�>�����w�V�H���|��].��'���Xwj}����3����"AS�)37J*u�38BqN�'c�X?&���Ig`i�ҋX����@�ڗe'=M�Z%�Ұv�~������]�!��r���4�$2p�8����WT�j
�I��w��,ਤ+;p	��F����U�D�>i�ל��K�Q���fd���Ig`iZ鎬����Y�V��#q![���>��Ig`iZ鎬����Y�V��#q̘�K>۟��Ig`iZ鎬����Y�V��#q�7��5��3r����=Y��_Q2�+�Y�3�+��m\'�C�,P�gD���g9Z鎬����Y�V��#qA/��? ��M��eNd�]�!���1����mrB�Z��g�mAx}��Mf���9���q���U�pzl��a�:��Y+Xf�B�>�9�ﻋ-���C�M��N��.W���ۗx>��OޘMf���9���q���U�pzl��a�DKj��=�B�>�9�ﻋ-������#έx��3����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h���[m���~������a����N���#t����n�~����p�@����9)����K�d���tn�u�$d�I�v`J��U����+=����7�>D�c�lQ@��~�
�KT\�mɍw�B�I:׷�F�20)�_SsJjvCn������Y�
���h$�7�R?�6��%]����	���a�P;m̳��\�B�6O�%� z����K�9y^6gVW���%@�~� ���I�����+����>�G0�?�I.M1�7�$�������zEK#�E��Ǵ\�"k�-1�	E�RpN&�2�C����}d�&ʛ}D_��Gɋ|5��N���5�r/1ހĮ�J�z�30��G�$,Ek���J�j��v�x��W"����UK�B�%��ό�;�LȫԷ�/^�\MGl�<���{��ZT��6|�� =��_�Z�G�a}Cfx��V$�wpxR���B��Q"}Hi���#2�}����[��Y-��J��׍���o�B��^�H��7TB�7a	�����Y�
��3��X1�'�3�$ �#^�Vn���.,&	M��0�d�Sd��_�a���n�|WC��0�O���ͪYQ��(V�0r�����K�9y^6gVW���%@�~� ���I�����+����>�G0�Y���ծǦ�3y
�*����zEK#�E��Ǵk�?H�$�IX[��O2<������ #M�)��u��`�|�&�#�E�d��������y��Ld_���1[���K��&�|�G�2I�wp(��C�712��}ǞK=<^��`Y�F�����I��#��
Mcu�T�M�ڤ [�f!�)�X�j(�� ����n�
_��q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r$����Gd"��U"�̩��k&Q��8�'��j^ҩ#��u1k�Z%ktg[���I\�wJ�G�����|�q<�_��s�֙���ƕ�*A�d�fWF0�M�J��@�WF;���.�P �0u��s$y���9����
�g�쎌�&���a�;�$y<޼e]]�q,�$X�刢0�]��	��M ?ؤ:�{��?�d���&�Q�.<�xN�[�����d(����I�ͭ[E~�ӵ(r7�l}�aB�g���B�
�I���^��*��O�t�!��6jV4�B��ٴ�� C�Q�+^�v�M�]�c۴l�&�j/vV_^{�^IN�f�w>{e�y{�הr�p�o27��e���im��1B"�A�`�=�ȭ^0E���^��0�$�ð��Tv��	�ʹ����?h���,��
��x(�i��/R�������	սL��$��ƹ���c�Xg�Yn��[_�����*�H`�~������w �I��!2,�4�+�-d��o�����x'=��O��(����<����+��!���8h��]$o8�(R�2�Ŋ�NE���5����A�>�xR�(V�RDFR7��U�z	��3�o�f���(�|�$��rÏ	�k�g�[�uQw�=+�����F�IQC`�%�l%zy�!jg�~m�Z��t�=Grh���?Zkܼ����Q�?������foȅ��k��4��s�S�,ii���5[��̔����'�u�X��@�v��~%BC�'y���xťwJ�G�����|�q<�_��s�֙`w7jH/g�3�G��+6Qk`e\����^�m�.4���2m�4�B��ٴm��ɅL�J)��e�O�{�h�� C���ŀK2���ƕo�����h4c�P�F~YEp1��t;��>��"���������X��1k��-��?O��xT�Z��5 
i�p]���#����k������CyC)ݼ�?E�~�#sv�RS�6���U��-|�v�LRu���$-��cLS��@�X+[%H����Ä�G�W8.+���W�dv��oTN!�������dҔ���Z��(��b=�i嬀֍�K�E�ө���x����8\l#�c�ۦ ���uN�;*�_��{M�бe���AP��=��;�n�dO�c����32��ӆo��*P�l$n�J[i���;��&͞d��M��V\�d	� 	qc�j�)Q��j8HQ��e�z�����,�W�B3���B[=cX�}��}v�_�j&��Ϻ�#Y��2�R�	��q'���y���4�CB��g��ۺ�D�͵SMI� y�r?�R�v~-}K�A�>�2�@w�?��?h��C���U�3�J~��k���k�[ݝ�B�W����k��)�-M
)#G�&���� d�":��p�T����pz��Ї��}I����#Q*b�6Ob���h+v҉����p�]ءVd|��()�T�~�k,9�? ��m�y���*>��$��� W�h�y��,-u��ƹ��t�d��`��'�BZ�-�a�Y�h�ݝ�B�W�ܴ����e.L*�d�,1X{���fz�}w�_c���\�+\�.��=YE��u��m�}�W-�W���E?��"�j��$�Lb�I�;�����k��\��@�u]�MP�T�%Σ��ĝ+����3J���|���s�44ȵ�B�B*��wj˻Z�zWz\ٿ�6�PG&XU��ѐaYR�B�\����K:C��<U_��s�֙f����h��y{�הr�R_ǌ� N��r*0��� F*,ƌN�jK�I�q������/f.������Ut�\��D��_:�!S�x�J�<�0|k4�Ż�&ǥ��a���F߸��S�Ȍ{ɝV�z����WN�d7!qzo_<�b"E��_'V��	��yO8S��%��3��J�:��n�&�E�aYR�B�\����K­[W�\M�_��s�֙]V�#9%���WN�d7!S�x�J�<�0|k4�@[�_zβr�v�������Q�^�� Fڱ���EC;�s�w{\�S�Ĕ�ZӞ�'�|,kW�F�����4�G�D�6(!rһpl�;�w����*H��M��FF�T	����$73���'���)Q��)���1
g�t�z�?�y)���t�%��	#�I�U�@B��rBWy03H��[.7|L����\c�;�^HUB����yt���w� �w(�
5��qD�KZ�����[�ƭM�R6�C1�f˾��S�d������m�I�_�k�8�ם��ɚ���ʈ�����)Hߋ,D���@�wR�� ������t^���\�}g��?`-ʂRcL�h�����WN�d79���'�!�'/2�%ͭ�=㜝�����E̒KV��	��y��Q�f<������E���YD�	��P�S�bN��E��锏��Z�� '����X,"�-��*1�#�;�����4�;��|B0F��#,k|2�Ω��!N�'�y�G