// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

module tstrom (addr, enab, q );
parameter LPM_FILE = "u1.hex";
input [7:0] addr;
input enab;
output [14:0] q;

  
asyn_rom_256x15 
// synopsys translate_off
           #(LPM_FILE)
// synopsys translate_on
      u1  (.Address(addr), .Q(q), .MemEnab(enab));

endmodule
