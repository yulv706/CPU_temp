��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-@���rahZ����*����Aڄ��[�k�|��ў��q����_�F��LF ��F9�>�^��M��7�m���<f#�}N9�h��/���b�%`F���\Zx�8��E��v�w��)?�� ! ,��e��~(l꼁��z��I._�O�
.�Zk�g�[��j�]�����8ɳ������F�A�xs̻��N��H^!�Kl�m�+�6��*��1�v����o�T
u�/%�O�"�F��� ��`p\x[���!�`�(i3W0�`��Ѣ�'t���/�!���c���"��z��"�����P��G�-�M��k�R��?xA4��^�y������9J�4Dvor0����.�q/�{<�x�fr��c�ZKY���#Ь�����Њ<s 2���ڠns6��������-VL�ސ���ƣ�L�/�\��9��IY���MTF�O;.��{C��|^����Yt��Z�M*q�M�/�-dOrS��E�����������I �x�r:�㜦��F?��߫�-H�/��� a�ik��Wʔ-�Y=.�"�K����X��֑xGV�M��T�t���(�zK�X饿��!��v����oX�$Z-�*��E��@��+'}���5M�YYroEێJR�VÀC�A��o��xȋ�l#ž��h�/,��ۿ����r�m�mIH3:Zt%��m&<�����9G�Ds|r�2?�����҃�F�� c��(�U�=��TA���#mԃw��+M}����j�����������d ���ѡ=�����Y �\Yy��V)�.�6C���Fz�k�좏1Y�_�R�|t�_=���$ۓ�����|Ǐ:�ues���$q��mKx"E&��� ��l$���D��Lh�Ԫ�u#7zǾIZ�Wl��>�;6W����F-P�u��.tƹy<c![���=$$h�8C& a�bD�G���O%���a\Y�����ḓ���X�,4�?n�[$��Q��3�O�2���Ė�� �Ueۡ萓'�al��p9�W�H{�G����g.Q�Q�?uG�)K|e�P4��&`��z��`5|⡰����r!�~WiZ��@Ő��thw��2r��h���\h��*�����g]��u�H1և���Bw��*`�|��K�z��}	�ʥ���S~:�:��3���C�P������eZ���(�Ow��/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@�ޗ9(����	�^��i���Ӿ���2���عf#�}N9�h�C����Y�q/L"t|Y�f�sJ�F���s�V�����<o�nïi�q{�f��a�:&�>��s���� T�8m��U}�	=�C��a���\�vūx`��:�r�^K������О.<�Ȭzn�w�'n�^0o����y�]��ӳ�Y�
Z�J
_�ʆ�In��tCF���y7�j�2\�{U�x���hA�4I^J<��H��&�ګvA���P`�|��K�zփZ���0�jݭ�F���h����tL���+��g�ڧZ��7�U�q��&�'n�^0of�`�(x���.j�,�3*������|���kJ_3#ڸZ鎬������rٮ�vF~�IK���Ig`i�ҋX����@�ڗe'���C1zh/�s��^a�T�~P�]k�!n}y���q���U�W����c�ZM�����{l�f|��rs�i�������k1T��v�܈�BT�^��a(􆿳�z��0������*�E��M@3%�w����$ĄҋX����`H���������h=-��;��lz������6�vg;Je'���Xw�j�7���|��{�r�\	��rR�^�V]��}R�wX�շ�R�������X��֑xGV�>�,2���7G#+�Ǘ0z�cUL�JJ�4(o�a\Y�����BT�^��a(􆿳��[ihC���%�ɏ�X,���֑xGV֚�X��M�TD���rs�i�>�Ca��?�o>�E]�٩��7�v�ԯ�`�L�i�C6�=�����!���;����J��6�vg;Je'���Xwb��Hg���'�r��'q�r.��c9�6�vg;Je'���Xw���e�KL[�#����KW�*�	S۱��J��q�P ڨ��S���Q�V�ɶ�w��V�k�j��ugM$BX���[��e��I�p\�WB�*�d��[� J���k�?�z7���%]��g���nU��X|Qeu��<�q{�f��a��\/�V����7�i���K�f�
�`�*%0�U�L�#_��^�+�J��;ۂ��IÙ=�HL'�kXyig@�����t��y�|�qx�]�V��v��K.Ū�C���D��j�69�$7��I[�x�]�V��v��K.Ū�C���D��^W�3B7��I[�x�]�V��v��K.Ū�C���DvW� �H`T7��I[�x�]�V��v��K.Ū�C���D�ӗ>���	7*6i��l!1�9���9M��I�� '����1��L��TZ����3;֍��@=;U�5V�˅|��k����z�KdL��[B�����؅��FJ��o�C���j��Ǌ�C��q�����/�~u+hBn�Y?v�<�!n}y��Y�{'%s�rOw������y$[|���"X��[z���6��+�x���+�qbp@���=ީa)��Ig`i�ҋX����f̲Az��%f�rE�X�e��Ig`i�ҋX����L$�����/���Ŋ�Ӑp�Dtq��Ig`i�ҋX����L$�����/���Ŋ��t��͝�u���Ig`i�ҋX����L$�����/���Ŋ����]D��;�č�Y���S�)37J*u�,�JL��ޅǐL�T�z�d6���|�_3#ڸZ鎬����Ĺ#{��	_1:Є8�Q;�m���!n}y��p�VU��Jm�QA�Q* �2��5���3(~s)tK��{l�f|��:2QYeƈ|���
p��v��֭��Ig`i�ҋX����L$�����/�Mv!���xl`�݃�|��].��'���Xw�����C�B�n}x��&�������{l�f|��:2QYeƈ�=�<�^\�c*�=|�WT�j
�I��w��,�,�JL���o:ϓ�gM��7P��T��TD���rs�i��ZIp����M�O��6a(􆿳� w�6p�d�H9M\��e���S��L�|[8�6�%ˮ�m�x���� ���S��S��6��o���+�@{fT�U�L�#_���29a���Q;5B5Y+�Y��d庒�D83��|��Yr���˩���.|�A6�E���?�.aݑMf���9���U� ���_j0��.@.�.H9���e#�|r�Mf���9���U� ���_j0��.@.�.H9���j��
�Mf���9���U� ���_j0��.@.�.H9��("�4��i�=�@��[�^������̇ki�D����m޴��eh�T�� �����r��T�,�'+���c[�u���褻��_j���=���a���Ѐ�uw�@.G5O7� ���Jg�C>��č�Y���S�)37J*uc�A�L'��-�S(�_Ma�~�Ǔ8���/�zeU�D�W�MԲ�����{l�f|�ό���.�܉��n* �w�-}�<��z��}�<ͧ�:|K5�w�x��?�����Ig`i�ҋX����L$�����/l◈�,��K.,�v�~������]�!���\B��V���)�xm���NX�c�|��].��'���Xw�����C����q
�o-x��az�d*�!n}y��p�VU��Jm�QA�Q* ���$þ�č�Y���S�)37J*u�,�JL��ޅǐL�T�z�_Flzk��_3#ڸZ鎬����Ĺ#{���0Q���ќבa��@IE�U����S8�	�Ms��3�˷���T�\ �������>�F����U���>$o?~�8r�k�K%*$�N�,�вԺL�9�d�e?��>ڃ(1����L�Y&
��L�>��ϣ'm�e��N(I:\����N��y]�u|�1��?��9O�������H��Y�{'%s�O��W��[�$��X�l�Lɼ�,0=]^	�&������%*$�N�,� :�:���H��߬���_;@�M�~��"����Y��ף��:����DZ���)i9%� MjC�9����T����X��֑xGV�}y���]D�]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/�Yum�IʝQ�`)��kѶ���� 7⸠z�V[���>(��+ �\Yy��x�@eӎ��'������;b&��E���L��v�я̛��q������ �4���q���U�pzl��a��Y&��Y����C1zhg�����g��=Y��_Q2�+�YɢX�B���y%�ɏ�X,���֑xGV�U�(f�Z��L�4?@�T�q���U��s��d�\Hq�o�d@-[�v:v�o���+���5���L����;j����>^���o���KEd��]^X0��
x-	���'�$HgL��)�J����f5i�A��I`��=J'����r
���I}}3M�C,����|#^�Vn����o[���=^��>D�c�lQ�����+�7끍J�[T�)��
�6���.�֌���<�a)�m�d�so�}a�C�ub;�;��V�k�j��ugM$BX;Ά\C��ɧ���7�)a���%}D�����!��g�-��\��OA�=�~�]��d�Y��o�6�֟�Zl��F�������WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zl��Ͳ�8�3���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂f#�}N9�h�C���ߠ���Y��EMܓ���;�e >���l�n�Zl��Ͳ�8�3
�{�-�>��t��ԱͽP�nT�N�+��9�M�s�F�:��8�^�.eO��q��S;gK�^~�U�'��gk=��[BfP3�e���b��M��Wv�'/B{�;4fx��V$�w�}MX�]y�Z��h��`�����o���c���w�L�R����*("ԛF�=���*� ��XLVt����G��5�On"WW��z&��y@���v���f��-/�J�¬��b����Lc�TH������7��ZΪm�T˚�Jz�0���je�Vmf��}S���u�����!�.3հjdo59
4/�]��	�`М��Wa;@��{�;F�~� �ne�Y�m�±��m|��Ѧ�#D�0[�H�l��}�Se[��[�$��X�l�Lɼ�:?-�2��$1&O����$ڭ�!�Mn�g�5'KL[����g_mWW�q1��MpM���Tf����Q1���bF���	i"�]/���я�40��YS�k�� �9*z@�o	�Au�����ώM:��2�n�ڤ���[U�&�n�.ZVRѿUJ�b��nw;�Z�/�k<����o��Ժ��e���S2x�FR���f5�%{ؕgD�%u?-/=z�ǀ��=�u���Fy�J~���;A���W�>����V;5h���X �8�4��Q>��~$�q����!��ZB^j��R��%T3��W< %�~3h���X ����C1zh/�s��^a�T�~P�]k��/h�Q-h���X ����X��֑xGV�96�O�n\�c*�=|�uFsY�w碪(���/��m�±��m|'�q�Om�@[�_zβr�v������t@���OHǙ <�E�t0��[y�Pm["QG�P�U��!�Mn�g�{�[>N�sr�S�
մtS5E]��:�L�������-VL��W�& :�L���R̶���[�σ8��i�	-_����l�Tc���v�I�	Zg� 1���XѤ�탎�Ŝ-���W	��X����' �Ϟ)kR��=��:�ݸ��~���W����@h~S܄= I>�-��}�x���5�DHb8��B�����̳9�o��j��")s
B�ݔ�]<�SIT������A��g��?qA��s��-��|a�,�)�*�.���3� 2dF.F?�o>�<���-,��V�F�P�_�^���\�}C6�=�����!���6�:�(�a�=�<�^�%&^�nƒg�|R��q� 8
�g��xsq��?�d���&�z��ܰ�S�P�s�a&�p�>��_5�L3�-bS�G�z8����?��0SߖP�s�a&�p�>��_5�L3�-bS����2F���|��{�r�\	��rR�,�o���,����Z�וzj7i�j��YoX���Q�ֱ�<�!5�k���������@%�:6ɬe�D�9N�j$���X��WG ���J
1�0�-��;���ݕ�
�o�y��Nկ����s��U;4�8�ߧ\����W �-g	�X��d��S�!g�d���z��R����0w�-��;����hJ�L��I/��\]��a-6�Dav���p�x��֑xGV�lᯆ�d�n��뾦�p�-a�D͢fU�9�׏�����MFi��|�3;c�<�%&^�nƒg�|R��qu�V�D/����<��ЕB;����v1a{J����b���\L���dL7A�k�6�Е�$8w|����X>j�V����������-��;���ݕ�
�o���z��V�7���N�ЕB;�����D���|0zC�N��z�5M�YYroE��t��ܠ�2�"q�䊒�G�����������4�~$���Vx�]�,qV��	��y ��f"���p���T������A�]�L���
QP�Tl$����Q>�^2�����Vc2�����Vc2�����Vc�C0�M���ҳ�$!nL^g	���lv7�H^%o�(ZH4~��2�����Vc2�����Vc2�����Vc⮆��`O|?,~��5Qo�n<�![��6�X�|K�mb�Xm[ �tf�u�c5���B�Zwqa�EuK��1�G�Qc�k]m��\��M���؈��k�;4���߫�����X��A���#���f��!���I0���t-���>*�+�n6+��c}Ex
:g��a��")�/K�ʕ�ˤSW�-��qs�VY�*R��=�9�3�j�c�Q�9�&�Q�z�וy�ǥJ��ѰǕ%�[.��j�D�EH<J�B@������_��]1�ڤbщ~��_�����XZ�i�Aum$&a:�P\�5"3�L����e���pJ�I4�[X+�������!d��]�%]�@�}w�,��~��@0ӸQ/�Z>�����^O�--�xS>e�c.E���و�FU�P�����X���ڿG��� �ʎ)������@��Kv1��l�^����D�I{GKg�!�4�yV�RDFR7��$�i3�a��b�âI���?Zkܼ��6�z�
^��1���K!<�v/�h��v����)F�Z�u6�������x����N	����|'Uʦ9��T�}���e�k�^o�e7+���߬<U��U �K]��z���Tr���
^��D'ڂ�+�;��;�;���Jq����*��=@r`y�pѲ�0)g�:jA�I;�śEN�.5snY��:H�T�f�3t ��	���DP�>>ompb-�<�vd�̪u��e�	}BEO�b=PGlcd�qS�?�E!^��@��1�@ �~)=��?�g�t�qy��YGzW{��o���2e��`p�K.o���n�ڿG��� ����׆�Tr�>b�L2�,Z�K6ԁcQ�w�;��л�yoZ�P/�����-VLt��(�"�6��j�_��ـ6�/�qW��G�� ��:	�����A�]\ң��;�v%��!�a\Y���������^�!�T�.�QCs">*�%�ɏ�X,���֑xGV�05 S�s�le�]0��&|��W&":@[�_zβrv���� g��?qA��s��-��S���Yp-�E��,@�,-ڥ��-St��I=:"p[94�.�a����h�g���ޔ�=:��}�$;��|Bͺ�L�A)�I*�?��m�±��m|,:e�)��.d�7~��ۣ�'�Aw���;e��J_���$�c��莨@g�p�7�Ͽ�K��G��#.�`���K�NG���m���߮�� e8�~��#`�k�(�5�T#%��ɬc��WN9q��N̆Ѿɪ�K���h+]��~}���3泂�3'�LD��-��r��M������q�X��E<.��,\ަ�It}�0�.�,���p�y��﹈�iZ��� CY�?�o>��	b[�q�*U*�������S,���J�X-����|.���=ީa)�!��ZB��M��7i�@�ZZl	�YI܁��[?��J���B�Ա?���q��cy�7�����3�!`�mL��1�G�Qc?KPبH��2���л�5Zbz�Z�x�r�m�d5�͐�-��;�� �T[�[P�E��6(�TKe�n510*���r�B�,{��I*�?��m�±��m|�_��$*-�Ps_*�GqW�w��fD���l׳d4��q���U�h+���dz��>�W2�����Vc2�����Vc2�����Vcl��w&� �na������b�4��"��W�'�Y���2�����Vc2�����Vc2�����Vc.�
͹U�1K�J{�T��C;�����u��0��K����y��@Ő��t'�������m�&(|dP�ݗ�}P�n:dL/U���j	��
#:��#~���5�f�y�X�p����O�Y��`�� ��$%�s�=�yx\o\w�����-VL(�sg��z�
! R�7��1�G�Qc�k]m���}���ݼ��1�G�Qc�Q�ޚ�꠹�h���VU�簦!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.��v'gn���1�/��+GkۯΔ��Ig~��
]yJْl��]�Bh#ґ�Dy��7a	��������W;5B5Y+� �i7�sp>����S �=�[T�)���}0�st&���\�vūx`��:�r�^K������О.|��	(���zL͊�q���g@b8�}O��t:(� �>u;YW���\�vś��X&`�KF2I��U�-��qs�VY���ܴ�&��'n�^0o���x�̗�����H��@Ő��t�����-VL1~�u�p���ӳ�Y�
�U�q��&�'n�^0o����SVc��ӳ�Y�
����.C� T2��zL͊�q����7y��"�j|~��A�!`�u�!j;5B5Y+��q	k���Ak�$����v7�'��O�q�Yz��"�ձ[%�U��Q�f�!�+��7P��T�<��z��}�צ:�)��-��7�Sc�Q��~�z��e�K����{l�f|����%Hlܾ�zx�8���#�!� k&oA�\ֆ-�֥�� ���Ig`i�ҋX����0�a1i~J�5�#(�@�%PX��n&oA�\ֆa��M(��E��jh�m!��ʧ�9�x�^4/��?Ev�~������]�!���R�qSe4�uS�4q�
��n��7��!n}y���q���U��֎)A=�s��]b_3#ڸZ鎬����8�������F�!���Fi����o_3#ڸZ鎬�������l�T�|�1��?���HEcx������]�!��	Ǹ�y85�:V�Fx��Wǖg3ȓ8���/��x���9D���o�Z�Xh�c�Q�j+�B��oy�{��vvfۛ��Q�]�_sC[k:!L)=���&�.�?GQ�.�� u�}��R�v�s�t��7v�(_4�Gé�ĻP�q����q�:��,��]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/��0��>d�0Q���g���C1zho)��
�ҋX������S8�^�8��nG�`�|��K�z&H�[&-n�g��U-�e�c����o0Q���g
3K������rg�D7�ҋX���� 
���u�ح(������O��X��M�TD���rs�i�>�Ca��?�o>�E]�٩��7�v�ԯ�`�L�iָt���(�x�_S1�����o�>�5��(�
t�������2�b]�iz�;Fuu�p�w4�i��������q�P ڨ��S���Q�V�ɶ�w���+GkۯΔ��Ig~��
]yJ�I�p\�WB������|q�谱O��\#+��SХ`�MϦ��pCeu��|��;ۂ���v8��j���	�$@ܫ�H9�&p�)����w&8��`Cq��p��=="vY0JߺGD@�F��qW��Ґ�Yj��2�+~c���<�"vY0JߺGD@�F��qW��Ґ�Yj��2�+~Ie��%�"vY0JߺGD@�F��qW��Ґ�Yj��2�+~m�����§���3;֍��@=;U�U�됵��D�oI��쬨L�|Hj����o��-�괂���I/���M��#�z�KdL��[B�����؅��FJ��o�C���j��Ǌ�C��q�����]����+g���wƱL<��z��}�0z�cULm�%������:F�X?�g��U-�e�4o��0��5K�������|��].��'���Xw����#�㬲C^�!n}y��p�VU��Jp��T����uD��^�3(~s)tK��{l�f|��:2QYeƈ|���
p�c�+�%I���Ig`i�ҋX����L$�����/l◈�,� Q���/v�~������]�!���\B��V���)�xmG�z"�!�_3#ڸZ鎬����Ĺ#{����$xN�In�(�At]�<��z��}�<ͧ�:|��u�읛���_H����č�Y���S�)37J*u�,�JL���o:ϓ�gM��7P��T��TD���rs�i��ZIp����M�O��6a(􆿳� w�6p�d�H9M\��e���S��%�e�J^}��A�"��ZbMHmH�ސ����6��o���+�@{fT�U�L�#_���29a���Q;5B5Y+�Y��d庒�D83��|��Yr���˩���.|�A6�E�@�,R����W�F��F�zL͊�q���19TH��M��oP�8��e�*��1�9���9M��C�0:���H����.���e홈t�T��1�9���9M��C�0:���H����:�(���i��t�T��1�9���9M��C�0:���H����y}�� ��t�T��1�9���9M��C�0 ��؋�[D����m޴��eh�T�� ������*ӶљvF�G�4�
Q`?�+G�	x��?,~x�]�V��v��K.Ū��)ZP1�^�=�Q��&9ʙ�~b��F�I5v�~������]�!��	Ǹ�y85���Vԓ4��[Ø�;�x�s�f޸��ބLȄ��'#�	��h�k�����p߷T�!n}y���q���U����G��e ݀�â�{l�f|��:2QYeƈ�WH���20��������e ݀�â�{l�f|��:2QYeƈ�WH���205�Gٙ��O�g�9��{l�f|��:2QYeƈ�WH���20��T��������Ia�i<��z��}�<ͧ�:|��u�읛Q)�2R}���č�Y���S�)37J*u�,�JL��ޅǐL�T�zʹ-j�b_3#ڸZ鎬����Ĺ#{���g�.���㱩� ���|��].��'���Xw�����C��m�U�I��W��!���{l�f|��:2QYeƈ�c�Z�~��i
E�v�~������]�!���\B��V���)�xm�0T���|��].��'���Xw�����U�\���P����^�i����(�
t��p�VU��Jm�QA�Q* 510*���8k>6s����]�!��	Ǹ�y85���Vԓ4��[Ø�;�x\�HP@�a����U�p��
���)��ZbMHmH�� �R�H��z���8�n��$���?\$��M��t9�<ݻ�\#+��SХ`�MϦ��pCeu��|��;ۂ���v8��j���	�$@ܫ�H9�&p�)����w&8��`Cq��p��=="vY0JߺGD@�F��qW��Ґ�Yj��2�+~c���<�"vY0JߺGD@�F��qW��Ґ�Yj��2�+~Ie��%�"vY0JߺGD@�F��qW��Ґ�Yj��2�+~@�����ϲ~X��t� ������ui���k ��؋�[D����m޴��eh�T�� ��������"
��xW�:R�yU�L�#_����Y7�Z�1�9���9M��C�0� 9��@f i#@���%&E����T�;��s\ڽ_3#ڸZ鎬�������(�����7$��t�Ȯ��ߊ���ł�!r��ބLȄ��'#�	��h�k�����p߷T�!n}y���q���U�>�(}%@��7�������{l�f|��:2QYeƈ�=�<�^��Q*J�<IjT%q�#�<��z��}�<ͧ�:|��ΥT�t֝��{�EG_3#ڸ�]�!���\B��V���)�xmB����B���|��].��'���Xw�����C�����d�W��!���{l�f|��:2QYeƈ�c�Z�~��i
E�v�~������]�!���\B��V���)�xm��B�ZE��|��].��'���Xw�����C�D> Υͤ���Ig`i7G#+�Ǘ0z�cULm�%������:F�X?�g��U-�e��!��'���GljJ��ƟWT�j
�I��w��,���|HH9M\��e���S���"
�	��d��4ɀ��ʶݦ�[:���BmIթ}bTm��0NB?��g��I��'�õ�Y���<�&4]��W[�f;q�sJHn��z�������a\Y�����|�i׋}%����v7Sx:����P�9�e�X�$Z-�*�����-VL}G�� �ܡ�)��nA6��>���pzl��a��8��*z�Sx�lޞ�ό���.�Q{�+�.�0]��;�A�f�A{XOl7}��G��C�C�.�.�\k�{j�$ bާ�kU�Mf���9���q���U�pzl��a������ґ�y�x��d~N�\'���Xw�2Qk�>	��6/z��\Ef�>��.���'���Xwa'�<� \E��T�ij���G��]_$Mf���9���q���U�KX�U~�?:h������BD|�	Sx�lޞ��rs�i�\_3�'����i� �߰a�P�Fpw��BT�^���8�B���z�C��йt�����,N���>S�`2dvϞ�]�!���1����m�n�\l�߅'O�%�3�ql��J�d�٣��5*���ӡ�.W���ۗ�5oMf���9���q���U�pzl��a��F��ţ<�Eg�N>Z9�8�4�X�'���Xwd�n]N�aB!�7a�0�:�5Ӡ�&H�[&-nD�P�E6���Qs��������(�=�ِmd��
/��y;���x/��\�d�٣�����6>���ZLl�]�z��"�����P��G�ޯ��ytaZ鎬����Y�V��#q5�31n�(?i˸3��Pư��]�!���1����m*�wX8�������p��~{pn˳T�ﻋ-���C�M��N��|�F7�_����'��e��"���N�@G�"Q��'���Xwa'�<� \%5�Ψa����g�cЉ�M��'ˑ�sO�rs�i�>�Ca��?�o>�E]�٩��7�v�ԯY��kB��d�o�P2}�).;��L�O#t����n��y,d��6{a�t P�^�\MGl�<���{��ZT��6|�� =��_�Z�G�a}Cfx��V$�w�Wή�li|��Q"}Hi���#2�}����[��Y-��J��׍���
�6���.�H��7TB�7a	�����Y�
��3��X1�'�3�$ �#^�Vn@j�cq9��M��0�d�Sd��_�a���n�|W���9IlcO���t���y1���?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��Le��	I���]�HЦ��EMW!���4m~�����c-�z��~��D:ǯ3�4���X�E��	�'�J���U�2Gޣסe� <���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9�xV��	7����G��O�L̍5��+'}����4L"�x��R�>(��F��eTQ�ȋ�V���w	����h _;��i�1�Q�^�� g�!�{5ܛ�	��A����¥��bMݪ��V�����׷eh��S�=�"�56RmHX���!���H���vO�[Jf퀔�������sr���0G3�,�ʗ2�Roܗw�m��%�۪�����s�x�9��喐Hj�Y�_�]	5�e� $p\�>���S�w҄�|5��s�#��v@���Jք�=�[��]�Kt�E*�#�,���ns)��E�$'/B{�;4{r�X��B&`��z��`?�d���&��W�!�ٱ��'��gk=���G��yʼ�	���Ek��d�/={ۀ�4����!oyY��&���t��@�����I���w�0\��.�gIt�!�����o����&�|�G�2�Ӑ�l���v����o��4��6�`!�A���
+,I�2Sj�	�$ɜ�\�۟�-?�d���&����{ԕ�h7�{`��������* -��ed.:E������ƄH����[��2����s�ZZ{�^�#�ZeT����7�@�0�r���a�)Z,�9�GKP�2�����Vc2�����Vc2�����Vcj+�;H,�^��Q��+I�[���ca��&�&-�(ZH4~��2�����Vc2�����Vc2�����VcSd�*-}Q��kL=�F>��o����o�fon�_�(�8�"�~;ѥ�RKW�*�	S^�����&s��חo���^hY'm0���?*е�^���wƄ�{Ƨ\bT]��7ۺ�#�����~��l��1aΉ����ߚ�����}�A,�S|��4���dq�e$��ӳ�Y�
ۼ��	K���$�(�+�G(��Y�Vd�8��N��(��{̑6ԉCy�8j�Y����I�k�%E~���J��ҝ���O�B���\媠 �eqɟ�R��(Q�u�<�w�i���2XC$2/G1�ԠֱTU8-R�T���k����$�����K�ֽ*�e��J-�1�q��)��b�Q�G��-�siË�M{z�(�˷�p"�.����L1�%Ŗ��g��T�/���B^�!n����d_��s����I8ԗx f�g\��*���?��c��R�?��Xq_í�F�s-w�?��?h�F�UΘ���.\��g(4��4�S�.u
i*�TWT0z��~�(E�POlb��]q������WV�#a�}!Z<>��V��&|6�łZ��0yI�[	ϱϭ����y>��v����jht��g�����9�g�klʟ���Q��:'�TPs_*�Gq�p���xg����6�������C;����Es���F1xk�k���L݁#g�k��g?	��o^3�|J�܄��� M{��(:/�b�&�q��ث#*�	���vAb@/��r �>/�w-���V��&|6�łZ��0yI�[	ϱ�f;[���v����jht��g��倉r˲���[yfX��[b%Ɨ�^Zp����4��x:A4b��JB䶓�([��}qn
V~$��|�;�#klʟ������u�h1�@/��r ��%�z�J����C���Uȓ�z�������C��R*E���&�Ut�\�8�8��gv8(?i˸3�J�
�MɂMv!���xP�o��x*ȩ��>d���,f1P�y�B���2L��x�ԉ�>B�R���>_�{�Z՟|
[;T�!'ؔsy1�n��뾦�f ;h�Z�O�#��K��%r]�Bа���/��D��c�Z�~c�}���Fo|k�LbB�R���>_c�Zਧ�%z��"�����P��G�Q"���_ނMv!���x8�8��gv8(?i˸3�J�
�M�'٥��gV�J�1���K���L���4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY�c���1�ā�����-ĭ5�6_ �nޝ3���� ��ɔ������?���;�$Y$E�B٘�#g�k��5د�������f�����X�G[ᱽәBe!^p��X��ئ,\ަ�It�_���U�L�#_���29a���Q������<`�y�����Cn%�}AU�L�#_��^�+�J����������@	Qg�m>�`^���t��˳�M:��2�;�琾BT���h�}q���'U�	�YI܁��DCX�.C��1�gB�� o� c �d�N9N�510*���IxoҢbu�g��A�i�8�=w��ir肃r���4�磕shf(�`�X�G[��c�fm���3�%Uo�'�D��¹��g�0�u
��"�!�sp�	O�ƻ��W\D�F3���%Ff"�	-7���ү��d�<��7���n���&�Pݭ��%�x �ǤZb�`�y�������"�X���G�����:�5Ӡ�X���e��
Ut�\�5�UI1�gB�� ]�Q%�n��뾦��"L?���P�o��x*ȩ��>d���,f1P�y�B���2L��\n0�8�:䩒=]'���76S=f�?TY�ސ�����)G�J�cbp��'@
9��y��%��3��ןmnRYpW����@	Q�M��k\z�$Y�G_Q#j<��#���z4�����i=���[taT��bX��WG ��v����jht��g��倉r˲���[yfX��[b%Ɨ�m��"���@��b_їE����ݾ-/���b練5د������
#>:����0^�� ŷ�[�}Gz�F:�@"��]����ڙ�����r(H\�ܢ��,	սL��$����,�ǰ���[�F/$�J���3Dm��A���%'ף'������d�l�'�al��paf��pD��>tT��N-بS� �D���B]���L�����=4�&��Q(I��M@3%�	����,�czb^y0�, bާ�kU��sC���X�45إ��ZWuȅ��SZ�N����VM�d�ꂕ0.p/��sH�}ˮіs�����������,hg~W#_pCeu��|̙1ږ���[�$��X�aM0��x9@xi�n��\ؤ�z;��$v��g�>�;6W�e�9�s[�A���t��˳.D,����	�YI܁��X����{o��&��;��L�Bza��i�g����l�1�ԀU�k�L�Z9@�;{�����%����%9��T�ِmd���u�a��bZ1�C�O�hh���X ��Y�����Y'b�'=�(�Ō����,��5si|�1��?�WdM4@�Z���}h
�#mԃw���k]m��yʥb�9ɮ2�����Vc2�����Vc2�����Vcv�iL�D��u]%_�ل�����5IΫN}q�~#�\��V2�����Vc2�����Vc2�����Vc.�
͹U�M�C:4�ֈґ�y�x�Q��C�uS�4q�
t�DY��b8!�ì�	jM�C:4���"r�V����U����r��<Н<�Xo���$����?�܃^�Y1V�&�i�д �rH:F��
 {�L_k6�iUrx���p#�r6�x5�A,I�@�"|VD.�+���s�f�I�w�U��|���1?�g��VĚ�d�>I�~�щ�X~��`O�g�q	G�Q��q�ﲾ�Bە��'��e����9�����Q�b6��pB0�iY�<�C7F�=j������<Va����7.N�ӃHF��v_}M������}'�=�+!�"y�W��n�)��o'>���?����u;϶i6����R�KL���:� #F�E�Zgu�t�1g��X��ن�	�a�B�����3����L�Y&Kfȵ3�\=�r}�Wq�ꑉ�� �3��l��gS#�-�tS~1x0PAok��G��]_$A�õ�٭�����ґ�y�x�l<Gt���{�]���q�GR��'Sդ�!��_S1�����o�>�5�Ǜ��k����>�lIorǟD�uiM���	�fmt����]$�﹈�i�~�Ԣ��D{5���U�L�#_��,Vit�-kݔ�yN{-v\L��"��#nS#y����m�(�����p߷Td��#���~$�q����!��ZB����=�+K�������үf�D r�f��h�3(~s)tK�h�RZ9�Y`�ِ{o�7���B�=�7�V���үf�D=�
�a�� D��ﺣ�i��¹ ^��y}$�)`� ��qQ��R��-���fx�Z�0�ԋ�Ƭ�����D�� >r�Z	�Ia���F�笣�.Z;�������xa��rװ� t��]�qa]�݊3�m�E;���20ӠH��=w�A2ޮ}'�=��~6��_��jt0��Ƅ^�=�]�_Jz������D��ܒ0�=1E�Êp!!v*!��4�b�Eƃ��Q-s�b!��u���͂EC�y��Q28U�sQ��=d�Ɇ�X�$Z-�*�����-VL�z����9�j��f6&��?N����Sr� �A����ҹ��)U��XI��ׅy&�Zz�IÛ	���~��s��>�̔���c�(�3��[��\*n6�-�Ƙw���+t�a���`������w�=u�A��7X_��7��W`i�X�QK6�E����*��[�$��X�l�Lɼ���C�O�d�xǬa��u����9A���q�O�����¯�P��C	,��Ȃ�	�����'C`ø�X�t�G�����u�����&�܁�^����r
��Cݮ2�����sE���y1+�줥G��j�D�EH<J�B@��(�hS�}e�܍ˢO�bF_��a��Mz���O?�Sկw��[#M�4�!�["[:����!��lSԃ�0�!𨱹�I*�?��m�±��m|�Mpl�p�;�s�*�:�L�������-VL�++��Lm�>�Q�k^�ïw��O�$Fg�#辭aE߅'O�%�z2�^4�l���lp����0�Rݯz"��G���P�f���oH�pNM�M��K�t0�5�]ؗ���0�E>�z�>C��?\$��M��ݺ|��W�_�\�Zr�2��_:��y$[|�h���X �õ�Y���<�&4]��W�q}�w|�/U���!-�iP��G��\OL^��>%�Нo@���;1?�[F�sp֟kh�y��;��lMԲ���L��S-�����$þh���X �����R]Y�3�#�����T<�t�S�@�l��tt�G�d�d�+��b2������ȼ�4�!O7I�"h#�)���w%e�D�m	$�WI��)A�
��v����=�\[L�R�X��Uq2��Z^��:�C�7�]���GljJ���a�X�� ��v|�ˑ����p|3�f0{��
�� �:&��L&fL0