-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.


--

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY TRIBUF_a8251 IS
    PORT (
        in1 : IN std_logic;
        oe  : IN std_logic;
        y   : OUT std_logic);
END TRIBUF_a8251;

ARCHITECTURE behavior OF TRIBUF_a8251 IS
BEGIN
    PROCESS (in1, oe)
    BEGIN
        IF oe'EVENT THEN
            IF oe = '0' THEN
                y <= TRANSPORT 'Z'  ;
            ELSIF oe = '1' THEN
                y <= TRANSPORT in1  ;
            END IF;
        ELSIF oe = '1' THEN
            y <= TRANSPORT in1  ;
        END IF;
    END PROCESS;
END behavior;

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DFF_a8251 IS
    PORT (
      	 d   : IN std_logic;
      	 clk : IN std_logic;
      	 clrn: IN std_logic;
      	 prn : IN std_logic;
      	 q   : OUT std_logic := '0');
END DFF_a8251;

ARCHITECTURE behavior OF DFF_a8251 IS
BEGIN

    PROCESS (clk, clrn, prn)
        VARIABLE result : std_logic := '0';
    BEGIN
        ASSERT NOT (prn = '0' AND clrn = '0')
            REPORT " prn and clrn both '0' on DFF"
            SEVERITY Warning;

        IF prn = '0' AND clrn = '1' THEN
            result := '1';
        ELSIF prn = '1' AND clrn = '0' THEN
            result := '0';
        ELSIF rising_edge(clk) THEN
            IF d = '1' OR d = '0' THEN
                result := d;
            END IF;
        END IF;

        IF result /= 'X' THEN
            q <= TRANSPORT result  ;
        END IF;

    END PROCESS;
END behavior;

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY FILTER_a8251 IS
    PORT (
        in1 : IN std_logic;
        y: OUT std_logic);
END FILTER_a8251;

ARCHITECTURE behavior OF FILTER_a8251 IS
BEGIN

    y <= in1;
END behavior;

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE work.tribuf_a8251;
USE work.dff_a8251;
USE work.filter_a8251;

ENTITY a8251 IS
    PORT (
      DIN : IN std_logic_vector(7 downto 0);
      DOUT : OUT std_logic_vector(7 downto 0);
      CLK : IN std_logic;
      CnD : IN std_logic;
      EXTSYNCD : IN std_logic;
      nCS : IN std_logic;
      nCTS : IN std_logic;
      nDSR : IN std_logic;
      nRD : IN std_logic;
      nRESET : IN std_logic;
      nRXC : IN std_logic;
      nTXC : IN std_logic;
      nWR : IN std_logic;
      RXD : IN std_logic;
      nDTR : OUT std_logic;
      nEN : OUT std_logic;
      nRTS : OUT std_logic;
      RXRDY : OUT std_logic;
      SYN_BRK : OUT std_logic;
      TXD : OUT std_logic;
      TXEMPTY : OUT std_logic;
      TXRDY : OUT std_logic);
END a8251;

ARCHITECTURE REVISION1_2 OF a8251 IS

SIGNAL gnd : std_logic := '0';
SIGNAL vcc : std_logic := '1';
SIGNAL
    n_83, n_84, n_85, n_86, n_87, a_G118_aOUT, n_89, n_90, n_91, n_92, n_93,
          n_94, a_G701_aOUT, n_96, n_97, n_98, n_99, n_100, n_101, a_G705_aOUT,
          n_103, n_104, n_105, n_106, n_107, n_108, a_G491_aOUT, n_110, n_111,
          n_112, n_113, n_114, n_115, a_G495_aOUT, n_117, n_118, n_119, n_120,
          n_121, n_122, a_G483_aOUT, n_124, n_125, n_126, n_127, n_128, n_129,
          a_G514_aOUT, n_131, n_132, n_133, n_134, n_135, n_136, a_G708_aOUT,
          n_138, n_139, n_140, n_141, n_142, n_143, a_STXRDY_aNOT_aQ, n_145,
          n_146, n_147, n_148, n_149, n_150, a_STXEMPTY_aNOT_aQ, n_152, n_153,
          n_154, n_155, n_156, n_157, a_STXD_aOUT, n_159, n_160, n_161, n_162,
          n_163, n_164, a_SSYN_BRK_aOUT, n_166, n_167, n_168, n_169, n_170,
          n_171, a_SRXRDY_aQ, n_173, n_174, n_175, n_176, n_177, n_178, a_SCMND_OUT_F5_G_aQ,
          n_180, n_181, n_182, n_183, n_184, n_185, a_SNEN_aNOT_aOUT, n_187,
          n_188, n_189, n_190, n_191, n_192, a_SCMND_OUT_F1_G_aQ, n_194, a_N580_aNOT_aOUT,
          a_N580_aNOT_aIN, n_197, n_198, n_199, a_N607_aOUT, n_201, a_LC1_C2_aOUT,
          n_203, a_SMODE_OUT_F3_G_aQ, a_SMODE_OUT_F3_G_aCLRN, a_SMODE_OUT_F3_G_aD,
          n_212, n_213, n_214, n_215, n_216, a_N82_aNOT_aOUT, n_218, a_N1034_aNOT_aOUT,
          n_220, n_221, n_222, a_SMODE_OUT_F3_G_aCLK, a_LC2_C16_aOUT, a_LC2_C16_aIN,
          n_227, n_228, n_229, a_N1189_aOUT, n_231, n_233, n_234, a_SMODE_OUT_F2_G_aQ,
          a_SMODE_OUT_F2_G_aCLRN, a_SMODE_OUT_F2_G_aD, n_242, n_243, n_244,
          n_245, n_246, n_247, n_248, n_249, n_250, n_251, a_SMODE_OUT_F2_G_aCLK,
          a_N1804_aQ, a_N1804_aCLRN, a_N1804_aD, n_260, n_261, n_262, a_N1807_aQ,
          n_264, n_265, a_N1804_aCLK, a_N1807_aCLRN, a_N1807_aD, n_273, n_274,
          n_275, n_277, n_279, n_281, n_282, a_N1807_aCLK, a_LC8_C7_aOUT,
          a_LC8_C7_aIN, n_286, n_287, n_288, a_LC1_C7_aNOT_aOUT, n_290, a_N1121_aNOT_aOUT,
          n_292, a_SCMND_OUT_F4_G_aQ, n_294, n_295, n_297, n_298, n_299, a_SCMND_OUT_F4_G_aCLRN,
          a_SCMND_OUT_F4_G_aD, n_306, n_307, n_308, n_309, n_310, n_311, a_SCMND_OUT_F4_G_aCLK,
          a_N101_aOUT, a_N101_aIN, n_315, n_316, n_317, a_N1757_aQ, n_319,
          a_N1756_aQ, n_321, a_N227_aNOT_aOUT, a_N227_aNOT_aIN, n_324, n_325,
          n_326, a_N130_aNOT_aOUT, n_328, a_N1165_aOUT, n_330, n_331, a_SMODE_OUT_F6_G_aQ,
          n_333, a_LC5_C20_aOUT, a_LC5_C20_aIN, n_336, n_337, n_338, a_N1754_aQ,
          n_340, n_341, n_342, n_343, n_344, n_345, n_346, a_N239_aOUT, a_N239_aIN,
          n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, a_SMODE_OUT_F7_G_aQ,
          n_358, n_359, a_N1754_aCLRN, a_N1754_aD, n_366, n_367, n_368, n_369,
          n_370, n_371, n_372, n_373, n_374, a_N1754_aCLK, a_N236_aOUT, a_N236_aIN,
          n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387,
          n_388, a_N1757_aCLRN, a_N1757_aD, n_395, n_396, n_397, n_398, n_399,
          n_400, n_401, n_402, a_N1757_aCLK, a_N235_aNOT_aOUT, a_N235_aNOT_aIN,
          n_406, n_407, n_408, n_409, n_410, n_411, n_412, a_N1756_aCLRN,
          a_N1756_aD, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426,
          n_427, n_428, a_N1756_aCLK, a_N1806_aQ, a_N1806_aCLRN, a_N1806_aD,
          n_437, n_438, n_439, a_N1808_aQ, n_441, n_442, a_N1806_aCLK, a_N1808_aCLRN,
          a_N1808_aD, n_450, n_451, n_452, mode_cmplt_aOUT, n_454, n_455,
          n_456, n_457, n_458, a_N1808_aCLK, a_N1898_aQ, a_N1898_aCLRN, a_N1898_aD,
          n_468, n_469, n_470, n_471, n_472, a_N1898_aCLK, a_N1897_aQ, a_N1897_aCLRN,
          a_N1897_aD, n_482, n_483, n_484, n_485, n_486, a_N1897_aCLK, a_N310_aNOT_aOUT,
          a_N310_aNOT_aIN, n_490, n_491, n_492, a_N296_aNOT_aOUT, n_494, a_SMODE_OUT_F0_G_aQ,
          n_496, n_497, n_498, a_SMODE_OUT_F1_G_aQ, n_500, a_LC3_B16_aOUT,
          a_LC3_B16_aIN, n_503, n_504, n_505, a_N1107_aOUT, n_507, a_N414_aQ,
          n_509, a_N413_aQ, n_511, n_512, a_N298_aOUT, n_514, n_515, n_516,
          a_N411_aQ, a_N411_aCLRN, a_N411_aD, n_524, n_525, n_526, a_N81_aNOT_aOUT,
          n_528, n_529, n_530, n_531, n_532, n_533, n_534, a_N411_aCLK, a_LC5_B18_aOUT,
          a_LC5_B18_aIN, n_539, n_540, n_541, a_N470_aOUT, n_543, a_N869_aQ,
          n_545, n_546, a_LC2_B11_aOUT, n_548, a_N606_aQ, n_550, a_N179_aOUT,
          a_N179_aIN, n_553, n_554, n_555, a_SSYNC2_F0_G_aQ, n_557, a_N729_aQ,
          n_559, n_560, n_561, a_SSYNC1_F0_G_aQ, n_563, a_N1093_aNOT_aOUT,
          a_N1093_aNOT_aIN, n_566, n_567, n_568, a_N1114_aNOT_aOUT, n_570,
          n_571, n_572, n_573, a_N2031_aQ, n_575, a_N869_aCLRN, a_N869_aD,
          n_582, n_583, n_584, n_585, a_N221_aNOT_aOUT, n_587, n_588, n_589,
          n_590, n_591, n_592, n_593, a_N869_aCLK, a_N1904_aQ, a_N1904_aCLRN,
          a_N1904_aD, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610,
          a_N1904_aCLK, a_N1903_aQ, a_N1903_aCLRN, a_N1903_aD, n_619, n_620,
          n_621, n_622, n_623, a_N1903_aCLK, a_LC6_C3_aOUT, a_LC6_C3_aIN,
          n_627, n_628, n_629, n_630, a_N1123_aNOT_aOUT, n_632, n_633, a_SMODE_OUT_F4_G_aQ,
          a_SMODE_OUT_F4_G_aCLRN, a_SMODE_OUT_F4_G_aD, n_641, n_642, n_643,
          n_644, n_645, n_646, n_647, n_648, n_649, n_650, a_SMODE_OUT_F4_G_aCLK,
          a_LC1_C3_aOUT, a_LC1_C3_aIN, n_654, n_655, n_656, n_657, n_658,
          n_659, n_661, a_SMODE_OUT_F6_G_aCLRN, a_SMODE_OUT_F6_G_aD, n_668,
          n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, a_SMODE_OUT_F6_G_aCLK,
          a_SCMND_OUT_F6_G_aQ, a_SCMND_OUT_F6_G_aCLRN, a_SCMND_OUT_F6_G_aD,
          n_686, n_687, n_688, n_689, a_N701_aNOT_aOUT, n_691, n_692, n_693,
          n_694, n_695, n_696, n_697, a_SCMND_OUT_F6_G_aCLK, a_N1895_aQ, a_N1895_aCLRN,
          a_N1895_aD, n_706, n_707, n_708, n_709, n_710, a_N1895_aCLK, a_N1811_aQ,
          a_N1811_aCLRN, a_N1811_aD, n_719, n_720, n_721, a_N1812_aQ, n_723,
          n_724, a_N1811_aCLK, a_N100_aOUT, a_N100_aIN, n_728, n_729, n_730,
          a_LC5_C13_aOUT, n_732, n_733, n_734, a_N1812_aCLRN, a_N1812_aD,
          n_741, n_742, n_743, n_744, n_745, n_747, n_748, n_749, a_N1812_aCLK,
          a_LC8_B20_aOUT, a_LC8_B20_aIN, n_753, n_754, n_755, n_756, n_757,
          a_SMODE_OUT_F5_G_aQ, n_759, n_760, n_761, n_762, n_763, n_764, n_765,
          n_766, n_767, n_768, n_769, n_770, n_771, a_LC4_B2_aOUT, a_LC4_B2_aIN,
          n_774, n_775, n_776, a_N1108_aNOT_aOUT, n_778, a_N1099_aNOT_aOUT,
          n_780, a_N1098_aNOT_aOUT, n_782, a_N1097_aNOT_aOUT, n_784, n_785,
          n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795,
          n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805,
          n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815,
          n_816, n_817, n_818, n_819, a_LC7_B2_aOUT, a_LC7_B2_aIN, n_822,
          n_823, n_824, a_N1096_aNOT_aOUT, n_826, a_N1095_aNOT_aOUT, n_828,
          a_N1094_aNOT_aOUT, n_830, n_831, n_832, n_833, n_834, n_835, n_836,
          n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846,
          n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856,
          n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866,
          a_N868_aQ, a_N868_aCLRN, a_N868_aD, n_874, n_875, n_876, n_877,
          n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887,
          a_N868_aCLK, a_LC5_B7_aOUT, a_LC5_B7_aIN, n_891, n_892, n_893, a_N1128_aNOT_aOUT,
          n_895, n_896, n_897, n_898, n_899, a_N616_aOUT, a_N616_aIN, n_902,
          n_903, n_904, a_LC8_B4_aNOT_aOUT, n_906, n_907, n_908, a_N80_aOUT,
          n_910, n_911, a_LC6_B7_aOUT, a_LC6_B7_aIN, n_914, n_915, n_916,
          a_N76_aNOT_aOUT, n_918, n_919, n_920, a_LC3_B7_aNOT_aOUT, n_922,
          a_LC8_B7_aOUT, a_LC8_B7_aIN, n_925, n_926, n_927, n_928, n_929,
          n_930, n_931, n_932, n_933, n_934, n_935, a_N414_aCLRN, a_N414_aD,
          n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951,
          n_952, a_N414_aCLK, a_LC2_B10_aOUT, a_LC2_B10_aIN, n_956, n_957,
          n_958, a_N1066_aNOT_aOUT, n_960, n_961, n_962, n_963, n_964, a_LC2_B4_aOUT,
          a_LC2_B4_aIN, n_967, n_968, n_969, a_N1179_aNOT_aOUT, n_971, a_N394_aQ,
          n_973, n_974, n_975, a_LC1_B4_aNOT_aOUT, n_977, n_978, n_979, n_980,
          a_N413_aCLRN, a_N413_aD, n_987, n_988, n_989, n_990, n_991, n_992,
          n_993, n_994, n_995, n_996, a_LC8_B10_aOUT, n_998, n_999, a_N413_aCLK,
          a_N1899_aQ, a_N1899_aCLRN, a_N1899_aD, n_1008, n_1009, n_1010, a_N1900_aQ,
          n_1012, n_1013, a_N1899_aCLK, a_N1900_aCLRN, a_N1900_aD, n_1021,
          n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, a_N1900_aCLK,
          a_SCMND_OUT_F0_G_aQ, a_SCMND_OUT_F0_G_aCLRN, a_SCMND_OUT_F0_G_aD,
          n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044,
          n_1045, n_1046, n_1047, a_SCMND_OUT_F0_G_aCLK, a_SRXREG_F0_G_aQ,
          a_SRXREG_F0_G_aCLRN, a_SRXREG_F0_G_aD, n_1056, n_1057, n_1058, a_N83_aOUT,
          n_1060, a_N79_aNOT_aOUT, n_1062, n_1063, n_1064, n_1065, a_N1100_aNOT_aOUT,
          n_1067, n_1068, n_1069, a_SRXREG_F0_G_aCLK, a_SRXREG_F1_G_aQ, a_SRXREG_F1_G_aCLRN,
          a_SRXREG_F1_G_aD, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083,
          n_1084, n_1085, a_N1101_aNOT_aOUT, n_1087, n_1088, n_1089, a_SRXREG_F1_G_aCLK,
          a_SRXREG_F2_G_aQ, a_SRXREG_F2_G_aCLRN, a_SRXREG_F2_G_aD, n_1098,
          n_1099, n_1100, n_1101, a_N134_aNOT_aOUT, n_1103, n_1104, n_1105,
          n_1106, a_N1102_aNOT_aOUT, n_1108, n_1109, n_1110, a_SRXREG_F2_G_aCLK,
          a_SRXREG_F3_G_aQ, a_SRXREG_F3_G_aCLRN, a_SRXREG_F3_G_aD, n_1119,
          n_1120, n_1121, n_1122, a_N1103_aNOT_aOUT, n_1124, n_1125, n_1126,
          n_1127, n_1128, n_1129, n_1130, a_SRXREG_F3_G_aCLK, a_LC7_A11_aOUT,
          a_LC7_A11_aIN, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, a_N1106_aNOT_aOUT,
          n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148,
          n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156,
          n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164,
          n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172,
          n_1173, n_1174, n_1175, n_1176, a_LC1_A11_aOUT, a_LC1_A11_aIN, n_1179,
          n_1180, n_1181, a_N1105_aNOT_aOUT, n_1183, n_1184, a_N96_aOUT, n_1186,
          n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194,
          n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202,
          n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210,
          n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218,
          n_1219, n_1220, n_1221, n_1222, a_N552_aNOT_aOUT, a_N552_aNOT_aIN,
          n_1225, n_1226, n_1227, a_N1104_aNOT_aOUT, n_1229, n_1230, n_1231,
          n_1232, n_1233, n_1234, a_N1998_aQ, n_1236, n_1237, n_1238, n_1239,
          n_1240, a_N551_aNOT_aOUT, a_N551_aNOT_aIN, n_1243, n_1244, n_1245,
          n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253,
          n_1254, n_1255, n_1256, a_LC2_C6_aOUT, a_LC2_C6_aIN, n_1259, n_1260,
          n_1261, n_1262, n_1263, n_1264, n_1265, a_LC5_C21_aOUT, a_LC5_C21_aIN,
          n_1268, n_1269, n_1270, n_1271, n_1272, pe_aQ, n_1274, n_1275, n_1276,
          n_1277, pe_aCLRN, pe_aD, n_1284, n_1285, n_1286, n_1287, n_1288,
          n_1289, n_1290, n_1291, n_1292, pe_aCLK, a_SRXREG_F4_G_aQ, a_SRXREG_F4_G_aCLRN,
          a_SRXREG_F4_G_aD, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306,
          n_1307, n_1308, n_1309, n_1310, n_1311, a_SRXREG_F4_G_aCLK, a_N325_aNOT_aOUT,
          a_N325_aNOT_aIN, n_1315, n_1316, n_1317, a_N1163_aNOT_aOUT, n_1319,
          a_N59_aQ, n_1321, a_N62_aQ, n_1323, a_N61_aQ, n_1325, n_1326, n_1327,
          n_1328, n_1329, a_N329_aNOT_aOUT, a_N329_aNOT_aIN, n_1332, n_1333,
          n_1334, a_N1183_aNOT_aOUT, n_1336, a_N1145_aOUT, n_1338, a_N64_aQ,
          n_1340, a_N63_aQ, n_1342, a_LC3_D3_aOUT, a_LC3_D3_aIN, n_1345, n_1346,
          n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, a_LC6_D4_aOUT,
          n_1355, n_1356, oe_aQ, oe_aCLRN, oe_aD, n_1364, n_1365, n_1366,
          n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374,
          oe_aCLK, a_LC4_D20_aOUT, a_LC4_D20_aIN, n_1378, n_1379, n_1380,
          n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, a_SRXREG_F5_G_aQ,
          a_SRXREG_F5_G_aCLRN, a_SRXREG_F5_G_aD, n_1395, n_1396, n_1397, n_1398,
          n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, a_SRXREG_F5_G_aCLK,
          a_N708_aNOT_aOUT, a_N708_aNOT_aIN, n_1409, n_1410, n_1411, n_1412,
          n_1413, n_1414, a_N707_aNOT_aOUT, a_N707_aNOT_aIN, n_1417, n_1418,
          n_1419, n_1420, n_1422, n_1423, n_1424, n_1425, a_N141_aNOT_aOUT,
          n_1427, n_1428, fe_aQ, fe_aCLRN, fe_aD, n_1436, n_1437, n_1438,
          n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, fe_aCLK, a_LC1_C6_aOUT,
          a_LC1_C6_aIN, n_1448, n_1449, n_1450, n_1451, n_1452, a_SRXREG_F6_G_aQ,
          a_SRXREG_F6_G_aCLRN, a_SRXREG_F6_G_aD, n_1460, n_1461, n_1462, n_1463,
          n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, a_SRXREG_F6_G_aCLK,
          a_SRXREG_F7_G_aQ, a_SRXREG_F7_G_aCLRN, a_SRXREG_F7_G_aD, n_1479,
          n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487,
          n_1488, n_1489, a_SRXREG_F7_G_aCLK, a_LC4_C7_aOUT, a_LC4_C7_aIN,
          n_1493, n_1494, n_1495, a_N1120_aNOT_aOUT, n_1497, n_1498, a_SCMND_OUT_F3_G_aQ,
          n_1500, n_1501, a_N613_aOUT, n_1503, n_1504, a_SCMND_OUT_F3_G_aCLRN,
          a_SCMND_OUT_F3_G_aD, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516,
          n_1517, n_1518, n_1519, n_1520, a_SCMND_OUT_F3_G_aCLK, a_LC2_C4_aOUT,
          a_LC2_C4_aIN, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530,
          a_SMODE_OUT_F0_G_aCLRN, a_SMODE_OUT_F0_G_aD, n_1537, n_1538, n_1539,
          n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, a_SMODE_OUT_F0_G_aCLK,
          a_LC6_C4_aOUT, a_LC6_C4_aIN, n_1550, n_1551, n_1552, n_1553, n_1554,
          n_1555, n_1557, a_SMODE_OUT_F1_G_aCLRN, a_SMODE_OUT_F1_G_aD, n_1564,
          n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572,
          n_1573, a_SMODE_OUT_F1_G_aCLK, a_SNEN_aNOT_aIN, n_1576, n_1577,
          n_1578, n_1579, n_1580, a_N1810_aQ, a_N1810_aCLRN, a_N1810_aD, n_1588,
          n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, a_N1810_aCLK, a_N1809_aQ,
          a_N1809_aCLRN, a_N1809_aD, n_1603, n_1604, n_1605, n_1606, n_1607,
          a_N1809_aCLK, a_N102_aOUT, a_N102_aIN, n_1611, n_1612, n_1613, n_1614,
          n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, a_N2010_aQ, a_N2010_aCLRN,
          a_N2010_aD, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, a_N655_aOUT,
          n_1635, n_1636, n_1637, n_1638, a_N2010_aCLK, a_STXRDY_aNOT_aCLRN,
          a_STXRDY_aNOT_aD, n_1647, n_1648, n_1649, n_1650, a_N77_aNOT_aOUT,
          n_1652, n_1653, n_1654, n_1655, a_N489_aNOT_aOUT, n_1657, n_1658,
          a_STXRDY_aNOT_aCLK, a_N534_aNOT_aOUT, a_N534_aNOT_aIN, n_1662, n_1663,
          n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, a_N1136_aNOT_aOUT,
          n_1672, n_1673, a_LC3_B14_aOUT, a_LC3_B14_aIN, n_1676, n_1677, n_1678,
          n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686,
          a_STXEMPTY_aNOT_aCLRN, a_STXEMPTY_aNOT_aD, n_1693, n_1694, n_1695,
          n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, a_STXEMPTY_aNOT_aCLK,
          a_SRXRDY_aCLRN, a_SRXRDY_aD, n_1710, n_1711, n_1712, n_1713, n_1714,
          n_1715, n_1716, n_1717, n_1718, n_1719, a_SRXRDY_aCLK, a_SCMND_OUT_F5_G_aCLRN,
          a_SCMND_OUT_F5_G_aD, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732,
          n_1733, n_1734, n_1735, n_1736, n_1737, a_SCMND_OUT_F5_G_aCLK, a_SCMND_OUT_F1_G_aCLRN,
          a_SCMND_OUT_F1_G_aD, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750,
          n_1751, n_1752, n_1753, n_1754, n_1755, a_SCMND_OUT_F1_G_aCLK, a_G118_aIN,
          n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765,
          n_1766, a_G701_aIN, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773,
          n_1774, n_1775, a_G705_aIN, n_1777, n_1778, n_1779, n_1780, n_1781,
          n_1782, n_1783, n_1784, a_G491_aIN, n_1786, n_1787, n_1788, n_1789,
          n_1790, n_1791, n_1792, n_1793, a_G495_aIN, n_1795, n_1796, n_1797,
          n_1798, n_1799, n_1800, n_1801, n_1802, a_G483_aIN, n_1804, n_1805,
          n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, a_SSYN_BRK_aIN,
          n_1813, n_1814, n_1815, a_N143_aOUT, n_1817, n_1818, n_1819, n_1820,
          n_1821, n_1822, n_1823, n_1824, n_1825, a_G514_aIN, n_1827, n_1828,
          n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, a_G708_aIN, n_1837,
          n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, a_N435_aOUT,
          a_N435_aIN, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853,
          n_1854, n_1855, n_1856, n_1857, a_N436_aOUT, a_N436_aIN, n_1860,
          n_1861, n_1862, n_1863, n_1864, n_1865, a_STXD_aIN, n_1867, n_1868,
          n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876,
          a_N1179_aNOT_aIN, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883,
          a_N76_aNOT_aIN, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890,
          a_N81_aNOT_aIN, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897,
          a_LC4_B6_aNOT_aOUT, a_LC4_B6_aNOT_aIN, n_1900, n_1901, n_1902, a_N365_aQ,
          n_1904, n_1905, a_N364_aQ, n_1907, a_LC7_B6_aNOT_aOUT, a_LC7_B6_aNOT_aIN,
          n_1910, n_1911, n_1912, a_N363_aQ, n_1914, n_1915, n_1916, a_LC3_B1_aNOT_aOUT,
          a_LC3_B1_aNOT_aIN, n_1919, n_1920, n_1921, a_N362_aQ, n_1923, n_1924,
          a_N360_aQ, n_1926, n_1927, n_1928, a_N361_aQ, n_1930, n_1931, n_1932,
          n_1933, n_1934, n_1935, n_1936, n_1937, a_N80_aIN, n_1939, n_1940,
          n_1941, a_N359_aQ, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948,
          n_1949, n_1950, a_N1136_aNOT_aIN, n_1952, n_1953, n_1954, n_1955,
          n_1956, n_1957, n_1958, n_1959, a_N470_aIN, n_1961, n_1962, n_1963,
          n_1964, n_1965, n_1966, a_LC3_B3_aOUT, a_LC3_B3_aIN, n_1969, n_1970,
          n_1971, n_1972, a_N599_aQ, n_1974, a_N311_aOUT, a_N311_aIN, n_1977,
          n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1985, a_N1064_aNOT_aOUT,
          a_N1064_aNOT_aIN, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993,
          n_1994, n_1995, a_LC1_B4_aNOT_aIN, n_1997, n_1998, n_1999, a_N396_aQ,
          n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, a_N397_aQ, n_2008,
          n_2009, n_2010, n_2011, n_2012, a_LC8_B4_aNOT_aIN, n_2014, n_2015,
          n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023,
          a_N1056_aOUT, a_N1056_aIN, n_2026, n_2027, n_2028, n_2029, n_2030,
          n_2031, n_2032, n_2033, a_N296_aNOT_aIN, n_2035, n_2036, n_2037,
          n_2038, n_2039, n_2040, n_2041, n_2042, a_N130_aNOT_aIN, n_2044,
          n_2045, n_2046, n_2047, n_2048, a_LC1_B8_aNOT_aOUT, a_LC1_B8_aNOT_aIN,
          n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058,
          a_N1114_aNOT_aIN, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065,
          n_2066, a_LC2_B7_aNOT_aOUT, a_LC2_B7_aNOT_aIN, n_2069, n_2070, n_2071,
          n_2072, n_2073, n_2074, n_2075, n_2076, a_LC3_B7_aNOT_aIN, n_2078,
          n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086,
          n_2087, a_N284_aOUT, a_N284_aIN, n_2090, n_2091, n_2092, n_2093,
          n_2094, n_2095, a_N1066_aNOT_aIN, n_2097, n_2098, n_2099, n_2100,
          n_2101, n_2102, n_2103, n_2104, a_N298_aIN, n_2106, n_2107, n_2108,
          n_2109, n_2110, n_2111, a_LC2_B16_aNOT_aOUT, a_LC2_B16_aNOT_aIN,
          n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121,
          a_LC5_B16_aNOT_aOUT, a_LC5_B16_aNOT_aIN, n_2124, n_2125, n_2126,
          n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134,
          n_2135, n_2136, n_2137, a_LC6_B1_aNOT_aOUT, a_LC6_B1_aNOT_aIN, n_2140,
          n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148,
          n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, a_LC4_B17_aNOT_aOUT,
          a_LC4_B17_aNOT_aIN, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163,
          n_2164, n_2165, n_2166, n_2167, n_2168, a_N1184_aNOT_aOUT, a_N1184_aNOT_aIN,
          n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, a_N1107_aIN, n_2178,
          n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186,
          n_2187, a_N1128_aNOT_aIN, n_2189, n_2190, n_2191, n_2192, n_2193,
          n_2194, a_N1065_aOUT, a_N1065_aIN, n_2197, n_2198, n_2199, n_2200,
          n_2201, n_2202, n_2203, n_2204, a_LC6_B16_aOUT, a_LC6_B16_aIN, n_2207,
          n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215,
          n_2216, a_N77_aNOT_aIN, n_2218, n_2219, n_2220, n_2221, n_2222,
          n_2223, n_2224, n_2225, a_N1032_aNOT_aOUT, a_N1032_aNOT_aIN, n_2228,
          n_2229, n_2230, n_2231, n_2232, n_2233, a_N221_aNOT_aIN, n_2235,
          n_2236, n_2237, n_2238, n_2239, a_N1134_aNOT_aOUT, a_N1134_aNOT_aIN,
          n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, a_LC5_C19_aOUT,
          a_LC5_C19_aIN, n_2250, n_2251, n_2252, n_2253, a_SSYNC1_F7_G_aQ,
          n_2255, n_2256, n_2257, n_2258, a_SSYNC2_F7_G_aQ, n_2260, n_2261,
          a_LC4_C19_aOUT, a_LC4_C19_aIN, n_2264, n_2265, n_2266, n_2267, n_2268,
          n_2269, n_2270, n_2271, n_2272, n_2273, a_N1138_aOUT, a_N1138_aIN,
          n_2276, n_2277, n_2278, n_2279, n_2280, a_N1108_aNOT_aIN, n_2282,
          n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, a_N2024_aQ,
          n_2291, a_N599_aCLRN, a_N599_aD, n_2298, n_2299, n_2300, n_2301,
          n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, a_N599_aCLK,
          a_LC2_B11_aIN, n_2311, n_2312, n_2313, n_2314, n_2315, a_LC4_B3_aOUT,
          a_LC4_B3_aIN, n_2318, n_2319, n_2320, n_2321, a_N601_aQ, n_2323,
          n_2324, n_2325, n_2326, a_LC3_C19_aOUT, a_LC3_C19_aIN, n_2329, n_2330,
          n_2331, a_SSYNC2_F6_G_aQ, n_2333, n_2334, n_2335, a_SSYNC1_F6_G_aQ,
          n_2337, n_2338, a_N1099_aNOT_aIN, n_2340, n_2341, n_2342, n_2343,
          a_N2025_aQ, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, a_N601_aCLRN,
          a_N601_aD, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363,
          n_2364, n_2365, n_2366, n_2367, a_N601_aCLK, a_LC5_B3_aOUT, a_LC5_B3_aIN,
          n_2371, n_2372, n_2373, n_2374, a_N602_aQ, n_2376, n_2377, n_2378,
          n_2379, a_N526_aOUT, a_N526_aIN, n_2382, n_2383, n_2384, n_2385,
          a_SSYNC1_F5_G_aQ, n_2387, n_2388, n_2389, n_2390, a_SSYNC2_F5_G_aQ,
          n_2392, n_2393, a_N1098_aNOT_aIN, n_2395, n_2396, n_2397, n_2398,
          n_2399, n_2400, n_2401, n_2402, a_N2026_aQ, n_2404, a_N602_aCLRN,
          a_N602_aD, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417,
          n_2418, n_2419, n_2420, n_2421, a_N602_aCLK, a_LC8_B2_aOUT, a_LC8_B2_aIN,
          n_2425, n_2426, n_2427, n_2428, a_N603_aQ, n_2430, n_2431, n_2432,
          n_2433, a_LC5_C18_aOUT, a_LC5_C18_aIN, n_2436, n_2437, n_2438, a_SSYNC2_F4_G_aQ,
          n_2440, n_2441, n_2442, a_SSYNC1_F4_G_aQ, n_2444, n_2445, a_N1097_aNOT_aIN,
          n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, a_N2027_aQ,
          n_2455, a_N603_aCLRN, a_N603_aD, n_2462, n_2463, n_2464, n_2465,
          n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, a_N603_aCLK,
          a_N1175_aNOT_aOUT, a_N1175_aNOT_aIN, n_2476, n_2477, n_2478, n_2479,
          n_2480, n_2481, a_N735_aNOT_aOUT, a_N735_aNOT_aIN, n_2484, n_2485,
          n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, a_LC5_D17_aOUT,
          a_LC5_D17_aIN, n_2494, n_2495, n_2496, a_N30_aQ, n_2498, n_2499,
          a_N28_aQ, n_2501, n_2502, n_2503, n_2504, a_N29_aQ, n_2506, n_2507,
          n_2508, n_2509, n_2510, n_2511, n_2512, a_N730_aNOT_aOUT, a_N730_aNOT_aIN,
          n_2515, n_2516, n_2517, a_N32_aQ, n_2519, n_2520, a_N31_aQ, n_2522,
          n_2523, a_N33_aQ, n_2525, n_2526, n_2527, a_LC2_D14_aOUT, a_LC2_D14_aIN,
          n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537,
          n_2538, n_2539, a_N83_aIN, n_2541, n_2542, n_2543, n_2544, n_2545,
          a_LC1_D14_aNOT_aOUT, a_LC1_D14_aNOT_aIN, n_2548, n_2549, n_2550,
          n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558,
          a_N1118_aNOT_aOUT, a_N1118_aNOT_aIN, n_2561, n_2562, n_2563, n_2564,
          n_2565, n_2566, a_N1149_aNOT_aOUT, a_N1149_aNOT_aIN, n_2569, n_2570,
          n_2571, n_2572, n_2573, n_2574, a_N89_aNOT_aOUT, a_N89_aNOT_aIN,
          n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584,
          a_N1163_aNOT_aIN, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591,
          a_N87_aNOT_aOUT, a_N87_aNOT_aIN, n_2594, n_2595, n_2596, n_2597,
          n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, a_N352_aOUT, a_N352_aIN,
          n_2606, n_2607, n_2608, n_2609, n_2610, a_N114_aOUT, a_N114_aIN,
          n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620,
          n_2621, n_2622, n_2623, a_N1144_aNOT_aOUT, a_N1144_aNOT_aIN, n_2626,
          n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634,
          n_2635, n_2636, n_2637, n_2638, n_2639, a_N95_aNOT_aOUT, a_N95_aNOT_aIN,
          n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, a_N155_aOUT, a_N155_aIN,
          n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657,
          n_2658, n_2659, a_LC2_D19_aOUT, a_LC2_D19_aIN, n_2662, n_2663, n_2664,
          n_2665, n_2666, n_2667, n_2668, n_2669, a_LC2_D17_aOUT, a_LC2_D17_aIN,
          n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679,
          n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687,
          a_LC5_D1_aOUT, a_LC5_D1_aIN, n_2690, n_2691, n_2692, n_2693, n_2694,
          n_2695, n_2696, n_2697, n_2698, n_2699, a_N116_aNOT_aOUT, a_N116_aNOT_aIN,
          n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709,
          n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, a_N751_aNOT_aOUT,
          a_N751_aNOT_aIN, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723,
          a_N1137_aNOT_aOUT, a_N1137_aNOT_aIN, n_2726, n_2727, n_2728, n_2729,
          n_2730, n_2731, a_LC4_D15_aOUT, a_LC4_D15_aIN, n_2734, n_2735, n_2736,
          n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, a_LC1_D15_aOUT,
          a_LC1_D15_aIN, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752,
          a_LC2_D15_aOUT, a_LC2_D15_aIN, n_2755, n_2756, n_2757, n_2758, n_2759,
          n_2760, n_2761, a_N1152_aNOT_aOUT, a_N1152_aNOT_aIN, n_2764, n_2765,
          n_2766, n_2767, n_2768, n_2769, a_LC5_D10_aOUT, a_LC5_D10_aIN, n_2772,
          n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780,
          n_2781, a_N1183_aNOT_aIN, n_2783, n_2784, n_2785, n_2786, n_2787,
          n_2788, a_N209_aOUT, a_N209_aIN, n_2791, n_2792, n_2793, n_2794,
          n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802,
          n_2803, n_2804, a_N207_aOUT, a_N207_aIN, n_2807, n_2808, n_2809,
          n_2810, n_2811, n_2812, a_N193_aNOT_aOUT, a_N193_aNOT_aIN, n_2815,
          n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, a_N153_aOUT,
          a_N153_aIN, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831,
          n_2832, n_2833, n_2834, a_N247_aNOT_aOUT, a_N247_aNOT_aIN, n_2837,
          n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, a_N743_aNOT_aOUT,
          a_N743_aNOT_aIN, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852,
          n_2853, n_2854, n_2855, n_2856, a_N125_aOUT, a_N125_aIN, n_2859,
          n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867,
          n_2868, n_2869, n_2870, n_2871, n_2872, a_N341_aOUT, a_N341_aIN,
          n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, a_N30_aCLRN,
          a_N30_aD, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894,
          n_2895, n_2896, n_2897, n_2898, a_N30_aCLK, a_N200_aOUT, a_N200_aIN,
          n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, a_N28_aCLRN, a_N28_aD,
          n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921,
          n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929,
          a_N28_aCLK, a_N29_aCLRN, a_N29_aD, n_2937, n_2938, n_2939, n_2940,
          n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948,
          n_2949, n_2950, n_2951, n_2952, a_N29_aCLK, a_LC5_B2_aOUT, a_LC5_B2_aIN,
          n_2956, n_2957, n_2958, n_2959, a_N604_aQ, n_2961, n_2962, n_2963,
          n_2964, a_LC5_C1_aOUT, a_LC5_C1_aIN, n_2967, n_2968, n_2969, a_SSYNC2_F3_G_aQ,
          n_2971, n_2972, n_2973, a_SSYNC1_F3_G_aQ, n_2975, n_2976, a_N1096_aNOT_aIN,
          n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, a_N2028_aQ,
          n_2986, a_N604_aCLRN, a_N604_aD, n_2993, n_2994, n_2995, n_2996,
          n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, a_N604_aCLK,
          a_N32_aCLRN, a_N32_aD, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016,
          n_3017, n_3018, n_3019, n_3020, n_3021, a_N32_aCLK, a_N31_aCLRN,
          a_N31_aD, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035,
          n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043,
          n_3044, a_N31_aCLK, a_N33_aCLRN, a_N33_aD, n_3052, n_3053, n_3054,
          n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062,
          a_N33_aCLK, a_N85_aNOT_aOUT, a_N85_aNOT_aIN, n_3066, n_3067, n_3068,
          n_3069, n_3070, n_3071, n_3072, n_3073, a_LC8_B10_aIN, n_3075, n_3076,
          n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084,
          n_3085, n_3086, n_3087, n_3088, a_N522_aNOT_aOUT, a_N522_aNOT_aIN,
          n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098,
          n_3099, n_3100, a_LC7_B10_aOUT, a_LC7_B10_aIN, n_3103, n_3104, n_3105,
          n_3106, n_3107, n_3108, n_3109, a_LC4_B10_aOUT, a_LC4_B10_aIN, n_3112,
          n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, a_LC1_B10_aOUT,
          a_LC1_B10_aIN, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127,
          n_3128, a_N365_aCLRN, a_N365_aD, n_3135, n_3136, n_3137, n_3138,
          n_3139, n_3140, n_3141, n_3142, n_3143, a_N365_aCLK, a_N364_aCLRN,
          a_N364_aD, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157,
          n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, a_N364_aCLK,
          a_N1189_aIN, n_3167, n_3168, n_3169, n_3170, n_3171, a_N82_aNOT_aIN,
          n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, a_N124_aOUT, a_N124_aIN,
          n_3181, n_3182, n_3183, n_3184, n_3185, a_N1035_aOUT, a_N1035_aIN,
          n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, a_LC1_C9_aOUT, a_LC1_C9_aIN,
          n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, a_SSYNC1_F5_G_aCLRN,
          a_SSYNC1_F5_G_aD, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214,
          n_3215, n_3216, n_3217, n_3218, a_SSYNC1_F5_G_aCLK, a_SSYNC1_F7_G_aCLRN,
          a_SSYNC1_F7_G_aD, n_3226, n_3227, n_3228, n_3229, n_3230, n_3232,
          n_3233, n_3234, n_3235, n_3236, n_3237, a_SSYNC1_F7_G_aCLK, a_LC2_C9_aOUT,
          a_LC2_C9_aIN, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247,
          a_SSYNC1_F6_G_aCLRN, a_SSYNC1_F6_G_aD, n_3254, n_3255, n_3256, n_3257,
          n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, a_SSYNC1_F6_G_aCLK,
          a_LC4_C9_aOUT, a_LC4_C9_aIN, n_3267, n_3268, n_3269, n_3270, n_3271,
          n_3272, n_3273, a_SSYNC1_F4_G_aCLRN, a_SSYNC1_F4_G_aD, n_3280, n_3281,
          n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289,
          a_SSYNC1_F4_G_aCLK, a_LC6_B18_aOUT, a_LC6_B18_aIN, n_3293, n_3294,
          n_3295, n_3296, a_N605_aQ, n_3298, n_3299, n_3300, n_3301, a_LC6_B19_aOUT,
          a_LC6_B19_aIN, n_3304, n_3305, n_3306, a_SSYNC2_F2_G_aQ, n_3308,
          n_3309, n_3310, a_SSYNC1_F2_G_aQ, n_3312, n_3313, a_N1095_aNOT_aIN,
          n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, a_N2029_aQ,
          n_3323, a_N605_aCLRN, a_N605_aD, n_3330, n_3331, n_3332, n_3333,
          n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, a_N605_aCLK,
          a_N129_aNOT_aOUT, a_N129_aNOT_aIN, n_3344, n_3345, n_3346, a_N919_aQ,
          n_3348, n_3349, n_3350, n_3351, a_N917_aQ, n_3353, n_3354, n_3355,
          n_3356, n_3357, n_3358, n_3359, n_3360, a_LC8_A9_aOUT, a_LC8_A9_aIN,
          n_3363, n_3364, n_3365, a_N920_aQ, n_3367, n_3368, a_N923_aQ, n_3370,
          n_3371, a_N921_aQ, n_3373, n_3374, a_N922_aQ, n_3376, a_N1126_aOUT,
          a_N1126_aIN, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385,
          n_3386, n_3387, n_3388, a_N919_aCLRN, a_N919_aD, n_3395, n_3396,
          n_3397, n_3398, n_3399, a_SCMND_OUT_F2_G_aQ, n_3401, n_3402, n_3403,
          n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411,
          a_N919_aCLK, a_N576_aOUT, a_N576_aIN, n_3415, n_3416, n_3417, n_3418,
          n_3419, n_3420, a_N564_aOUT, a_N564_aIN, n_3423, n_3424, n_3425,
          n_3426, n_3427, n_3428, n_3429, a_N1083_aOUT, a_N1083_aIN, n_3432,
          n_3433, n_3434, n_3435, n_3436, n_3437, a_N917_aCLRN, a_N917_aD,
          n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451,
          n_3452, n_3453, n_3454, n_3455, n_3456, a_N917_aCLK, a_LC5_A9_aOUT,
          a_LC5_A9_aIN, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, a_LC6_A9_aOUT,
          a_LC6_A9_aIN, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474,
          n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, a_N920_aCLRN, a_N920_aD,
          n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, a_N920_aCLK, a_N923_aCLRN,
          a_N923_aD, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506,
          n_3507, n_3508, n_3509, n_3510, a_N923_aCLK, a_N921_aCLRN, a_N921_aD,
          n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525,
          n_3526, n_3527, n_3528, a_N921_aCLK, a_N922_aCLRN, a_N922_aD, n_3536,
          n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544,
          n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, a_N922_aCLK,
          a_N489_aNOT_aIN, n_3554, n_3555, n_3556, n_3557, n_3558, a_N1197_aOUT,
          a_N1197_aIN, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, a_N1198_aOUT,
          a_N1198_aIN, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, a_N2027_aCLRN,
          a_N2027_aD, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587,
          n_3588, n_3589, a_N2027_aCLK, a_N2026_aCLRN, a_N2026_aD, n_3597,
          n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605,
          a_N2026_aCLK, a_N2025_aCLRN, a_N2025_aD, n_3613, n_3614, n_3615,
          n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623,
          a_N2025_aCLK, a_N2024_aCLRN, a_N2024_aD, n_3631, n_3632, n_3633,
          n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641,
          a_N2024_aCLK, a_N1165_aIN, n_3644, n_3645, n_3646, n_3647, n_3648,
          a_N608_aOUT, a_N608_aIN, n_3651, n_3652, n_3653, n_3654, n_3655,
          a_LC5_B5_aOUT, a_LC5_B5_aIN, n_3658, n_3659, n_3660, n_3661, n_3662,
          n_3663, a_N120_aOUT, a_N120_aIN, n_3666, n_3667, n_3668, n_3669,
          n_3670, a_SSYNC1_F1_G_aQ, a_SSYNC1_F1_G_aCLRN, a_SSYNC1_F1_G_aD,
          n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685,
          n_3686, a_SSYNC1_F1_G_aCLK, a_N1168_aNOT_aOUT, a_N1168_aNOT_aIN,
          n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, a_N1116_aNOT_aOUT,
          a_N1116_aNOT_aIN, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703,
          a_N718_aOUT, a_N718_aIN, n_3706, n_3707, n_3708, n_3709, n_3710,
          n_3711, a_SSYNC2_F1_G_aQ, a_SSYNC2_F1_G_aCLRN, a_SSYNC2_F1_G_aD,
          n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726,
          n_3727, n_3728, a_SSYNC2_F1_G_aCLK, a_N723_aOUT, a_N723_aIN, n_3732,
          n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, a_SSYNC2_F2_G_aCLRN,
          a_SSYNC2_F2_G_aD, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750,
          n_3751, n_3752, n_3753, n_3754, a_SSYNC2_F2_G_aCLK, a_N103_aOUT,
          a_N103_aIN, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, a_SSYNC1_F2_G_aCLRN,
          a_SSYNC1_F2_G_aD, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775,
          n_3776, n_3777, n_3778, a_SSYNC1_F2_G_aCLK, a_LC4_C5_aOUT, a_LC4_C5_aIN,
          n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, a_SSYNC2_F3_G_aCLRN,
          a_SSYNC2_F3_G_aD, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799,
          n_3800, n_3801, n_3802, n_3803, a_SSYNC2_F3_G_aCLK, a_N607_aIN,
          n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, a_SSYNC1_F3_G_aCLRN,
          a_SSYNC1_F3_G_aD, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824,
          n_3825, n_3826, n_3827, a_SSYNC1_F3_G_aCLK, a_N363_aCLRN, a_N363_aD,
          n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842,
          n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, a_N363_aCLK, a_N362_aCLRN,
          a_N362_aD, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862,
          n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, a_N362_aCLK,
          a_LC8_B1_aOUT, a_LC8_B1_aIN, n_3873, n_3874, n_3875, n_3876, n_3877,
          n_3878, a_N360_aCLRN, a_N360_aD, n_3885, n_3886, n_3887, n_3888,
          n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896,
          n_3897, n_3898, a_N360_aCLK, a_LC7_B1_aOUT, a_LC7_B1_aIN, n_3902,
          n_3903, n_3904, n_3905, n_3906, a_N361_aCLRN, a_N361_aD, n_3913,
          n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921,
          n_3922, n_3923, n_3924, n_3925, n_3926, a_N361_aCLK, a_N234_aNOT_aOUT,
          a_N234_aNOT_aIN, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935,
          n_3936, a_SSYNC2_F6_G_aCLRN, a_SSYNC2_F6_G_aD, n_3943, n_3944, n_3945,
          n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, a_SSYNC2_F6_G_aCLK,
          a_SSYNC2_F7_G_aCLRN, a_SSYNC2_F7_G_aD, n_3959, n_3960, n_3961, n_3962,
          n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, a_SSYNC2_F7_G_aCLK,
          a_N233_aNOT_aOUT, a_N233_aNOT_aIN, n_3973, n_3974, n_3975, n_3976,
          n_3977, n_3978, n_3979, a_SSYNC2_F5_G_aCLRN, a_SSYNC2_F5_G_aD, n_3986,
          n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994,
          a_SSYNC2_F5_G_aCLK, a_SSYNC2_F4_G_aCLRN, a_SSYNC2_F4_G_aD, n_4002,
          n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010,
          n_4011, n_4012, a_SSYNC2_F4_G_aCLK, a_N1120_aNOT_aIN, n_4015, n_4016,
          n_4017, a_N1902_aQ, n_4019, n_4020, a_N1901_aQ, n_4022, a_N1052_aOUT,
          a_N1052_aIN, n_4025, n_4026, n_4027, n_4028, n_4029, a_N1177_aOUT,
          a_N1177_aIN, n_4032, n_4033, n_4034, a_N1555_aQ, n_4036, a_N1556_aQ,
          n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, a_N420_aOUT, a_N420_aIN,
          n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053,
          n_4054, n_4055, a_LC3_A1_aOUT, a_LC3_A1_aIN, n_4058, n_4059, n_4060,
          n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068,
          n_4069, a_LC4_A1_aOUT, a_LC4_A1_aIN, n_4072, n_4073, n_4074, n_4075,
          n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083,
          a_N1050_aOUT, a_N1050_aIN, n_4086, n_4087, n_4088, n_4089, n_4090,
          n_4091, a_N1187_aOUT, a_N1187_aIN, n_4094, n_4095, n_4096, n_4097,
          n_4098, a_LC1_A15_aOUT, a_LC1_A15_aIN, n_4101, n_4102, n_4103, n_4104,
          n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112,
          a_N676_aOUT, a_N676_aIN, n_4115, n_4116, n_4117, n_4118, n_4119,
          n_4120, n_4121, n_4122, n_4123, n_4124, a_N1135_aNOT_aOUT, a_N1135_aNOT_aIN,
          n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, a_LC2_A15_aNOT_aOUT,
          a_LC2_A15_aNOT_aIN, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140,
          n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148,
          a_N425_aNOT_aOUT, a_N425_aNOT_aIN, n_4151, n_4152, n_4153, n_4154,
          n_4155, n_4156, n_4157, n_4158, n_4159, a_N1054_aNOT_aOUT, a_N1054_aNOT_aIN,
          n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169,
          a_N1049_aNOT_aOUT, a_N1049_aNOT_aIN, n_4172, n_4173, n_4174, n_4175,
          n_4176, n_4177, n_4178, n_4179, a_LC2_A1_aNOT_aOUT, a_LC2_A1_aNOT_aIN,
          n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, a_LC5_A1_aOUT, a_LC5_A1_aIN,
          n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197,
          a_N427_aOUT, a_N427_aIN, n_4200, n_4201, n_4202, n_4203, a_N1170_aQ,
          n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212,
          n_4213, n_4214, n_4215, n_4216, a_N423_aNOT_aOUT, a_N423_aNOT_aIN,
          n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, a_N428_aOUT,
          a_N428_aIN, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234,
          n_4235, n_4236, a_LC2_A12_aOUT, a_LC2_A12_aIN, n_4239, n_4240, n_4241,
          n_4242, a_N1169_aQ, n_4244, n_4245, n_4246, a_N1167_aQ, n_4248,
          n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, a_N132_aOUT, a_N132_aIN,
          n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, a_N1171_aQ, n_4264,
          n_4265, n_4266, n_4267, n_4268, n_4269, a_N1146_aOUT, a_N1146_aIN,
          n_4272, n_4273, n_4274, n_4275, n_4276, a_LC1_D2_aNOT_aOUT, a_LC1_D2_aNOT_aIN,
          n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286,
          a_N1070_aOUT, a_N1070_aIN, n_4289, n_4290, n_4291, n_4292, n_4293,
          n_4294, n_4295, a_LC5_C13_aIN, n_4297, n_4298, n_4299, n_4300, n_4301,
          n_4302, n_4303, n_4304, n_4305, n_4306, a_N127_aOUT, a_N127_aIN,
          n_4309, n_4310, n_4311, n_4312, n_4313, a_N1073_aNOT_aOUT, a_N1073_aNOT_aIN,
          n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323,
          n_4324, n_4325, a_N1072_aNOT_aOUT, a_N1072_aNOT_aIN, n_4328, n_4329,
          n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337,
          a_N1164_aOUT, a_N1164_aIN, n_4340, n_4341, n_4342, n_4343, n_4344,
          a_N1080_aOUT, a_N1080_aIN, n_4347, n_4348, n_4349, n_4350, n_4351,
          n_4352, a_LC5_D16_aOUT, a_LC5_D16_aIN, n_4355, n_4356, n_4357, n_4358,
          n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, a_N167_aOUT, a_N167_aIN,
          n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, a_N35_aNOT_aOUT,
          a_N35_aNOT_aIN, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381,
          n_4382, n_4383, a_N465_aNOT_aOUT, a_N465_aNOT_aIN, n_4386, n_4387,
          n_4388, n_4389, a_N1302_aQ, n_4391, n_4392, n_4393, a_N1301_aQ,
          n_4395, a_N1051_aOUT, a_N1051_aIN, n_4398, n_4399, n_4400, n_4401,
          n_4402, n_4403, a_N466_aNOT_aOUT, a_N466_aNOT_aIN, n_4406, n_4407,
          n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, a_N1303_aQ, n_4415,
          n_4416, n_4417, n_4418, a_N54_aOUT, a_N54_aIN, n_4421, n_4422, n_4423,
          n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, a_N12_aOUT,
          a_N12_aIN, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439,
          a_N1304_aQ, n_4441, n_4442, n_4443, a_N1102_aNOT_aIN, n_4445, n_4446,
          n_4447, n_4448, a_N1305_aQ, n_4450, n_4451, n_4452, n_4453, a_N1205_aOUT,
          a_N1205_aIN, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462,
          n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470,
          n_4471, n_4472, n_4473, a_N1_aOUT, a_N1_aIN, n_4476, n_4477, n_4478,
          n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, a_N456_aNOT_aOUT,
          a_N456_aNOT_aIN, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493,
          n_4494, n_4495, n_4496, n_4497, a_LC4_A11_aOUT, a_LC4_A11_aIN, n_4500,
          n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508,
          n_4509, a_LC3_A11_aOUT, a_LC3_A11_aIN, n_4512, n_4513, n_4514, n_4515,
          n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, a_LC4_A21_aOUT,
          a_LC4_A21_aIN, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4530,
          n_4531, a_N1306_aQ, n_4533, n_4534, a_N1101_aNOT_aIN, n_4536, n_4537,
          n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545,
          a_N145_aNOT_aOUT, a_N145_aNOT_aIN, n_4548, n_4549, n_4550, n_4551,
          n_4552, a_N161_aOUT, a_N161_aIN, n_4555, n_4556, n_4557, n_4558,
          n_4559, n_4560, n_4561, n_4562, a_LC5_A2_aOUT, a_LC5_A2_aIN, n_4565,
          n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573,
          n_4574, a_LC1_A21_aOUT, a_LC1_A21_aIN, n_4577, n_4578, n_4579, n_4580,
          a_N1307_aQ, n_4582, n_4583, n_4584, n_4585, a_LC5_A21_aOUT, a_LC5_A21_aIN,
          n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595,
          a_LC2_A21_aOUT, a_LC2_A21_aIN, n_4598, n_4599, n_4600, n_4601, n_4602,
          n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, a_N1100_aNOT_aIN,
          n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618,
          a_N1203_aOUT, a_N1203_aIN, n_4621, n_4622, n_4623, n_4624, n_4625,
          n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633,
          n_4634, n_4635, n_4636, n_4637, n_4638, a_LC4_B9_aNOT_aOUT, a_LC4_B9_aNOT_aIN,
          n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648,
          n_4649, n_4650, n_4651, n_4652, a_LC2_A10_aOUT, a_LC2_A10_aIN, n_4655,
          n_4656, n_4657, n_4658, n_4659, n_4660, a_N1300_aQ, n_4662, n_4663,
          a_N1039_aNOT_aOUT, a_N1039_aNOT_aIN, n_4666, n_4667, n_4668, n_4669,
          n_4670, n_4671, a_N398_aOUT, a_N398_aIN, n_4674, n_4675, n_4676,
          n_4677, n_4678, n_4679, n_4680, n_4681, a_LC6_A4_aOUT, a_LC6_A4_aIN,
          n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691,
          n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, a_N1040_aNOT_aOUT,
          a_N1040_aNOT_aIN, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705,
          n_4706, a_N687_aNOT_aOUT, a_N687_aNOT_aIN, n_4709, n_4710, n_4711,
          n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719,
          a_N1041_aNOT_aOUT, a_N1041_aNOT_aIN, n_4722, n_4723, n_4724, n_4725,
          n_4726, n_4727, a_N1105_aNOT_aIN, n_4729, n_4730, n_4731, n_4732,
          n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, a_N144_aNOT_aOUT,
          a_N144_aNOT_aIN, n_4742, n_4743, n_4744, n_4745, n_4746, a_N165_aOUT,
          a_N165_aIN, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755,
          n_4756, a_LC5_C12_aNOT_aOUT, a_LC5_C12_aNOT_aIN, n_4759, n_4760,
          n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768,
          n_4769, n_4770, n_4771, n_4772, a_N461_aNOT_aOUT, a_N461_aNOT_aIN,
          n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782,
          n_4783, n_4784, n_4785, n_4786, a_N458_aNOT_aOUT, a_N458_aNOT_aIN,
          n_4789, n_4790, n_4791, n_4792, n_4793, a_N22_aNOT_aOUT, a_N22_aNOT_aIN,
          n_4796, n_4797, n_4798, n_4799, n_4800, n_4801, a_N20_aNOT_aOUT,
          a_N20_aNOT_aIN, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809,
          n_4810, n_4811, n_4812, n_4813, a_N19_aNOT_aOUT, a_N19_aNOT_aIN,
          n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823,
          a_N55_aNOT_aOUT, a_N55_aNOT_aIN, n_4826, n_4827, n_4828, n_4829,
          n_4830, n_4831, n_4832, n_4833, a_N56_aNOT_aOUT, a_N56_aNOT_aIN,
          n_4836, n_4837, n_4838, n_4839, n_4840, a_N1103_aNOT_aIN, n_4842,
          n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850,
          n_4851, n_4852, a_N1206_aOUT, a_N1206_aIN, n_4855, n_4856, n_4857,
          n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865,
          n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, a_N96_aIN,
          n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, a_N166_aOUT, a_N166_aIN,
          n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889,
          a_LC2_C11_aNOT_aOUT, a_LC2_C11_aNOT_aIN, n_4892, n_4893, n_4894,
          n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902,
          n_4903, n_4904, n_4905, a_LC3_A19_aOUT, a_LC3_A19_aIN, n_4908, n_4909,
          n_4910, n_4911, n_4912, n_4913, a_LC1_A19_aOUT, a_LC1_A19_aIN, n_4916,
          n_4917, n_4918, n_4919, n_4920, n_4921, a_N1106_aNOT_aIN, n_4923,
          n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931,
          n_4932, n_4933, a_N686_aOUT, a_N686_aIN, n_4936, n_4937, n_4938,
          n_4939, n_4940, n_4941, n_4942, n_4943, a_N1077_aOUT, a_N1077_aIN,
          n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953,
          n_4954, n_4955, n_4956, n_4957, a_N694_aNOT_aOUT, a_N694_aNOT_aIN,
          n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967,
          a_N696_aNOT_aOUT, a_N696_aNOT_aIN, n_4970, n_4971, n_4972, n_4973,
          n_4974, n_4975, n_4976, n_4977, a_LC6_A19_aOUT, a_LC6_A19_aIN, n_4980,
          n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988,
          n_4989, a_N1104_aNOT_aIN, n_4991, n_4992, n_4993, n_4994, n_4995,
          n_4996, n_4997, n_4998, n_4999, n_5000, a_N1207_aOUT, a_N1207_aIN,
          n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010,
          n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018,
          n_5019, n_5020, a_N135_aOUT, a_N135_aIN, n_5023, n_5024, n_5025,
          n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, a_N1038_aNOT_aOUT,
          a_N1038_aNOT_aIN, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040,
          n_5041, n_5042, a_N1212_aOUT, a_N1212_aIN, n_5045, n_5046, n_5047,
          n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055,
          n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, a_N1210_aOUT,
          a_N1210_aIN, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071,
          n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079,
          n_5080, n_5081, n_5082, a_LC2_B9_aOUT, a_LC2_B9_aIN, n_5085, n_5086,
          n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094,
          n_5095, n_5096, a_LC1_C12_aOUT, a_LC1_C12_aIN, n_5099, n_5100, n_5101,
          n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109,
          n_5110, n_5111, n_5112, a_N1213_aOUT, a_N1213_aIN, n_5115, n_5116,
          n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124,
          n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132,
          a_LC1_C11_aOUT, a_LC1_C11_aIN, n_5135, n_5136, n_5137, n_5138, n_5139,
          n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147,
          n_5148, a_N1215_aOUT, a_N1215_aIN, n_5151, n_5152, n_5153, n_5154,
          n_5155, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162,
          a_N1214_aOUT, a_N1214_aIN, n_5165, n_5166, n_5167, n_5168, n_5169,
          n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177,
          n_5178, n_5179, n_5180, n_5181, n_5182, a_N1194_aNOT_aOUT, a_N1194_aNOT_aIN,
          n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192,
          n_5193, n_5194, a_N1037_aNOT_aOUT, a_N1037_aNOT_aIN, n_5197, n_5198,
          n_5199, n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, n_5206,
          a_LC6_A15_aOUT, a_LC6_A15_aIN, n_5209, n_5210, n_5211, n_5212, n_5213,
          n_5214, n_5215, n_5216, n_5217, a_N1125_aOUT, a_N1125_aIN, n_5220,
          n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228,
          n_5229, n_5230, a_N86_aOUT, a_N86_aIN, n_5233, n_5234, n_5235, n_5236,
          n_5237, n_5238, n_5239, a_N91_aOUT, a_N91_aIN, n_5242, n_5243, n_5244,
          n_5245, n_5246, a_LC8_D21_aOUT, a_LC8_D21_aIN, n_5249, n_5250, n_5251,
          n_5252, n_5253, n_5254, a_LC2_D7_aOUT, a_LC2_D7_aIN, n_5257, n_5258,
          n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, a_N524_aOUT, a_N524_aIN,
          n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274,
          n_5275, n_5276, n_5277, a_N1124_aNOT_aOUT, a_N1124_aNOT_aIN, n_5280,
          n_5281, n_5282, n_5283, n_5284, n_5285, a_N1170_aCLRN, a_N1170_aD,
          n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299,
          n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307,
          a_N1170_aCLK, a_N376_aOUT, a_N376_aIN, n_5311, n_5312, n_5313, n_5314,
          n_5315, n_5316, a_N1169_aCLRN, a_N1169_aD, n_5323, n_5324, n_5325,
          n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333,
          a_N1169_aCLK, a_N1167_aCLRN, a_N1167_aD, n_5341, n_5342, n_5343,
          n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351,
          n_5352, n_5353, n_5354, n_5355, n_5356, a_N1167_aCLK, a_N720_aOUT,
          a_N720_aIN, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365, n_5366,
          a_SSYNC2_F0_G_aCLRN, a_SSYNC2_F0_G_aD, n_5373, n_5374, n_5375, n_5376,
          n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, a_SSYNC2_F0_G_aCLK,
          a_N729_aCLRN, a_N729_aD, n_5390, n_5391, n_5392, n_5393, n_5394,
          n_5395, n_5396, n_5397, n_5398, n_5399, n_5400, n_5401, n_5402,
          a_N729_aCLK, a_N119_aOUT, a_N119_aIN, n_5406, n_5407, n_5408, n_5409,
          n_5410, a_SSYNC1_F0_G_aCLRN, a_SSYNC1_F0_G_aD, n_5417, n_5418, n_5419,
          n_5420, n_5421, n_5422, n_5423, n_5424, n_5425, a_SSYNC1_F0_G_aCLK,
          a_N2030_aQ, a_N2030_aCLRN, a_N2030_aD, n_5434, n_5435, n_5436, n_5437,
          n_5438, n_5439, n_5440, n_5441, n_5442, a_N2030_aCLK, a_N2029_aCLRN,
          a_N2029_aD, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456,
          n_5457, n_5458, a_N2029_aCLK, a_N2028_aCLRN, a_N2028_aD, n_5466,
          n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473, n_5474,
          a_N2028_aCLK, a_LC2_B1_aOUT, a_LC2_B1_aIN, n_5478, n_5479, n_5480,
          n_5481, n_5482, n_5483, n_5484, a_N359_aCLRN, a_N359_aD, n_5491,
          n_5492, n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499,
          n_5500, n_5501, n_5502, n_5503, n_5504, a_N359_aCLK, a_N396_aCLRN,
          a_N396_aD, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, n_5518,
          n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526,
          n_5527, a_N396_aCLK, a_N397_aCLRN, a_N397_aD, n_5535, n_5536, n_5537,
          n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545,
          a_N397_aCLK, a_N1171_aCLRN, a_N1171_aD, n_5553, n_5554, n_5555,
          n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562, n_5563,
          a_N1171_aCLK, a_LC3_A3_aOUT, a_LC3_A3_aIN, n_5567, n_5568, n_5569,
          a_N1553_aQ, n_5571, n_5572, n_5573, a_LC3_D4_aNOT_aOUT, a_LC3_D4_aNOT_aIN,
          n_5576, n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, a_LC4_D4_aOUT,
          a_LC4_D4_aIN, n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, a_LC2_D4_aOUT,
          a_LC2_D4_aIN, n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599,
          a_LC5_D4_aOUT, a_LC5_D4_aIN, n_5602, n_5603, n_5604, n_5605, n_5606,
          n_5607, n_5608, a_LC6_D4_aIN, n_5610, n_5611, n_5612, n_5613, n_5614,
          n_5615, n_5616, n_5617, n_5618, n_5619, a_N1145_aIN, n_5621, n_5622,
          n_5623, n_5624, n_5625, n_5626, a_N467_aNOT_aOUT, a_N467_aNOT_aIN,
          n_5629, n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636,
          n_5637, n_5638, n_5639, a_N113_aNOT_aOUT, a_N113_aNOT_aIN, n_5642,
          n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649, a_N79_aNOT_aIN,
          n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, a_LC2_A3_aOUT, a_LC2_A3_aIN,
          n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5665, n_5666,
          a_N1160_aOUT, a_N1160_aIN, n_5669, n_5670, n_5671, n_5672, n_5673,
          a_N1117_aOUT, a_N1117_aIN, n_5676, n_5677, n_5678, n_5679, n_5680,
          a_LC6_A3_aOUT, a_LC6_A3_aIN, n_5683, n_5684, n_5685, n_5686, n_5687,
          n_5688, a_N1553_aCLRN, a_N1553_aD, n_5695, n_5696, n_5697, n_5698,
          n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705, a_N1553_aCLK,
          a_N1307_aCLRN, a_N1307_aD, n_5713, n_5714, n_5715, n_5716, n_5717,
          n_5718, n_5719, n_5720, n_5721, n_5722, n_5723, a_N1307_aCLK, a_N1306_aCLRN,
          a_N1306_aD, n_5731, n_5732, n_5733, n_5734, n_5735, n_5736, n_5737,
          n_5738, n_5739, n_5740, n_5741, a_N1306_aCLK, a_N1069_aOUT, a_N1069_aIN,
          n_5745, n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, a_N59_aCLRN,
          a_N59_aD, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764,
          n_5765, n_5766, n_5767, n_5768, n_5769, a_N59_aCLK, a_N1302_aCLRN,
          a_N1302_aD, n_5777, n_5778, n_5779, n_5780, n_5781, n_5782, n_5783,
          n_5784, n_5785, n_5786, n_5787, a_N1302_aCLK, a_LC4_B18_aOUT, a_LC4_B18_aIN,
          n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798,
          a_N178_aOUT, a_N178_aIN, n_5801, n_5802, n_5803, n_5804, n_5805,
          n_5806, n_5807, n_5808, a_N1094_aNOT_aIN, n_5810, n_5811, n_5812,
          n_5813, n_5814, n_5815, n_5816, n_5817, a_N606_aCLRN, a_N606_aD,
          n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831,
          n_5832, n_5833, n_5834, a_N606_aCLK, a_LC4_A7_aOUT, a_LC4_A7_aIN,
          n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845,
          n_5846, n_5847, n_5848, a_LC2_A7_aOUT, a_LC2_A7_aIN, n_5851, n_5852,
          n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860,
          a_N134_aNOT_aIN, n_5862, n_5863, n_5864, n_5865, n_5866, a_N1193_aOUT,
          a_N1193_aIN, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874, a_N278_aOUT,
          a_N278_aIN, n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883,
          n_5884, n_5885, a_LC6_A13_aOUT, a_LC6_A13_aIN, n_5888, n_5889, n_5890,
          n_5891, n_5892, n_5893, a_LC2_A13_aOUT, a_LC2_A13_aIN, n_5896, n_5897,
          n_5898, n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905,
          a_N264_aNOT_aOUT, a_N264_aNOT_aIN, n_5908, n_5909, n_5910, n_5911,
          n_5912, n_5913, n_5914, n_5915, n_5916, n_5917, a_N1555_aCLRN, a_N1555_aD,
          n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931,
          n_5932, n_5933, n_5934, a_N1555_aCLK, a_LC4_A3_aOUT, a_LC4_A3_aIN,
          n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944, n_5945,
          a_LC5_A3_aOUT, a_LC5_A3_aIN, n_5948, n_5949, n_5950, n_5951, n_5952,
          n_5953, n_5954, n_5955, a_LC1_A3_aOUT, a_LC1_A3_aIN, n_5958, n_5959,
          n_5960, n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967,
          n_5968, a_LC5_A7_aOUT, a_LC5_A7_aIN, n_5971, n_5972, n_5973, n_5974,
          n_5975, n_5976, n_5977, a_N1556_aCLRN, a_N1556_aD, n_5984, n_5985,
          n_5986, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993,
          n_5994, a_N1556_aCLK, a_LC6_D13_aOUT, a_LC6_D13_aIN, n_5998, n_5999,
          n_6000, n_6001, n_6002, n_6003, a_N108_aNOT_aOUT, a_N108_aNOT_aIN,
          n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012, n_6013,
          mode_cmplt_aIN, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020,
          n_6021, a_LC6_D11_aOUT, a_LC6_D11_aIN, n_6025, n_6026, n_6027, n_6028,
          n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, a_LC5_D11_aOUT,
          a_LC5_D11_aIN, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043,
          n_6044, n_6045, a_LC7_D11_aOUT, a_LC7_D11_aIN, n_6048, n_6049, n_6050,
          n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, a_LC7_D10_aOUT,
          a_LC7_D10_aIN, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065,
          n_6066, a_LC4_D8_aOUT, a_LC4_D8_aIN, n_6069, n_6070, n_6071, n_6072,
          n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, a_N1158_aOUT, a_N1158_aIN,
          n_6081, n_6082, n_6083, n_6084, n_6085, a_N745_aNOT_aOUT, a_N745_aNOT_aIN,
          n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095,
          n_6096, n_6097, n_6098, a_LC3_D8_aOUT, a_LC3_D8_aIN, n_6101, n_6102,
          n_6103, n_6104, n_6105, n_6106, n_6107, n_6108, n_6109, n_6110,
          a_LC7_D7_aOUT, a_LC7_D7_aIN, n_6113, n_6114, n_6115, n_6116, n_6117,
          n_6118, a_N141_aNOT_aIN, n_6120, n_6121, n_6122, n_6123, n_6124,
          n_6125, n_6126, a_N106_aNOT_aOUT, a_N106_aNOT_aIN, n_6129, n_6130,
          n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, a_LC4_D10_aOUT,
          a_LC4_D10_aIN, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146,
          n_6147, n_6148, n_6149, a_LC5_D13_aOUT, a_LC5_D13_aIN, n_6152, n_6153,
          n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160, n_6161,
          a_N740_aNOT_aOUT, a_N740_aNOT_aIN, n_6164, n_6165, n_6166, n_6167,
          n_6168, n_6169, a_N64_aCLRN, a_N64_aD, n_6176, n_6177, n_6178, n_6179,
          n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, a_N64_aCLK, a_N1301_aCLRN,
          a_N1301_aD, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199,
          n_6200, n_6201, n_6202, n_6203, a_N1301_aCLK, a_N1998_aCLRN, a_N1998_aD,
          n_6211, n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6218,
          n_6219, n_6220, n_6221, a_N1998_aCLK, a_N1300_aCLRN, a_N1300_aD,
          n_6229, n_6230, n_6231, n_6232, n_6233, n_6234, n_6235, n_6236,
          n_6237, n_6238, n_6239, a_N1300_aCLK, a_N2031_aCLRN, a_N2031_aD,
          n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254,
          n_6255, a_N2031_aCLK, a_N1123_aNOT_aIN, n_6258, n_6259, n_6260,
          n_6261, n_6262, n_6263, n_6264, n_6265, a_LC3_C8_aOUT, a_LC3_C8_aIN,
          n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, a_N1034_aNOT_aIN,
          n_6276, n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283,
          a_SMODE_OUT_F5_G_aCLRN, a_SMODE_OUT_F5_G_aD, n_6290, n_6291, n_6292,
          n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, a_SMODE_OUT_F5_G_aCLK,
          a_N317_aOUT, a_N317_aIN, n_6303, n_6304, n_6305, n_6306, n_6307,
          a_N394_aCLRN, a_N394_aD, n_6314, n_6315, n_6316, n_6317, n_6318,
          n_6319, n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326,
          n_6327, n_6328, n_6329, a_N394_aCLK, a_N1067_aOUT, a_N1067_aIN,
          n_6333, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339, a_LC3_D10_aOUT,
          a_LC3_D10_aIN, n_6342, n_6343, n_6344, n_6345, n_6346, n_6347, n_6348,
          n_6349, n_6350, n_6351, a_LC2_D13_aOUT, a_LC2_D13_aIN, n_6354, n_6355,
          n_6356, n_6357, n_6358, n_6359, n_6360, n_6361, n_6362, a_LC4_D13_aOUT,
          a_LC4_D13_aIN, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371,
          n_6372, n_6373, a_N62_aCLRN, a_N62_aD, n_6380, n_6381, n_6382, n_6383,
          n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, a_N62_aCLK, a_LC1_C7_aNOT_aIN,
          n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, a_N1121_aNOT_aIN,
          n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, a_N701_aNOT_aIN,
          n_6407, n_6408, n_6409, n_6410, n_6411, a_N611_aOUT, a_N611_aIN,
          n_6414, n_6415, n_6416, n_6417, n_6418, a_N613_aIN, n_6420, n_6421,
          n_6422, n_6423, n_6424, n_6425, n_6426, n_6427, n_6428, n_6429,
          a_SCMND_OUT_F7_G_aQ, a_SCMND_OUT_F7_G_aCLRN, a_SCMND_OUT_F7_G_aD,
          n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443, n_6444,
          n_6445, n_6446, a_SCMND_OUT_F7_G_aCLK, a_N1902_aCLRN, a_N1902_aD,
          n_6454, n_6455, n_6456, n_6457, n_6458, a_N1902_aCLK, a_N1901_aCLRN,
          a_N1901_aD, n_6466, n_6467, n_6468, n_6469, n_6470, a_N1901_aCLK,
          a_N1305_aCLRN, a_N1305_aD, n_6478, n_6479, n_6480, n_6481, n_6482,
          n_6483, n_6484, n_6485, n_6486, n_6487, n_6488, a_N1305_aCLK, a_N1304_aCLRN,
          a_N1304_aD, n_6496, n_6497, n_6498, n_6499, n_6500, n_6501, n_6502,
          n_6503, n_6504, n_6505, n_6506, a_N1304_aCLK, a_N1303_aCLRN, a_N1303_aD,
          n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520, n_6521,
          n_6522, n_6523, n_6524, a_N1303_aCLK, a_LC3_C3_aOUT, a_LC3_C3_aIN,
          n_6528, n_6529, n_6530, n_6531, n_6532, n_6533, a_SMODE_OUT_F7_G_aCLRN,
          a_SMODE_OUT_F7_G_aD, n_6540, n_6541, n_6542, n_6543, n_6544, n_6545,
          n_6546, n_6547, n_6548, n_6549, a_SMODE_OUT_F7_G_aCLK, a_LC1_A8_aOUT,
          a_LC1_A8_aIN, n_6553, n_6554, n_6555, a_N965_aQ, n_6557, n_6558,
          a_N963_aQ, n_6560, n_6561, a_N964_aQ, n_6563, n_6564, a_N962_aQ,
          n_6566, a_LC4_A8_aOUT, a_LC4_A8_aIN, n_6569, n_6570, n_6571, n_6572,
          n_6573, n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, a_LC3_A8_aOUT,
          a_LC3_A8_aIN, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588,
          n_6589, n_6590, n_6591, n_6592, n_6593, n_6594, n_6595, a_N383_aOUT,
          a_N383_aIN, n_6598, n_6599, n_6600, n_6601, n_6602, n_6603, n_6604,
          n_6605, n_6606, n_6607, a_LC2_A8_aOUT, a_LC2_A8_aIN, n_6610, n_6611,
          n_6612, n_6613, n_6614, n_6615, n_6616, n_6617, n_6618, n_6619,
          n_6620, n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6627,
          n_6628, n_6629, n_6630, a_N390_aOUT, a_N390_aIN, n_6633, n_6634,
          n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641, n_6642,
          a_N143_aIN, n_6644, n_6645, n_6646, n_6647, n_6648, n_6649, n_6650,
          n_6651, n_6652, n_6653, n_6654, a_LC1_A6_aOUT, a_LC1_A6_aIN, n_6657,
          n_6658, n_6659, n_6660, n_6661, a_N451_aOUT, a_N451_aIN, n_6664,
          n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, a_N965_aCLRN,
          a_N965_aD, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684,
          n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692,
          n_6693, a_N965_aCLK, a_N455_aNOT_aOUT, a_N455_aNOT_aIN, n_6697,
          n_6698, n_6699, n_6700, n_6701, n_6702, a_N450_aOUT, a_N450_aIN,
          n_6705, n_6706, n_6707, n_6708, n_6709, a_N963_aCLRN, a_N963_aD,
          n_6716, n_6717, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723,
          n_6724, n_6725, n_6726, n_6727, n_6728, a_N963_aCLK, a_N964_aCLRN,
          a_N964_aD, n_6736, n_6737, n_6738, n_6739, n_6740, n_6741, n_6742,
          n_6743, n_6744, n_6745, n_6746, n_6747, n_6748, a_N964_aCLK, a_N962_aCLRN,
          a_N962_aD, n_6756, n_6757, n_6758, n_6759, n_6760, n_6761, n_6762,
          n_6763, n_6764, n_6765, n_6766, n_6767, n_6768, n_6769, n_6770,
          n_6771, a_N962_aCLK, a_LC7_C15_aOUT, a_LC7_C15_aIN, n_6775, n_6776,
          n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783, a_SCMND_OUT_F2_G_aCLRN,
          a_SCMND_OUT_F2_G_aD, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795,
          n_6796, n_6797, n_6798, n_6799, a_SCMND_OUT_F2_G_aCLK, a_N659_aNOT_aOUT,
          a_N659_aNOT_aIN, n_6803, n_6804, n_6805, n_6806, n_6807, n_6808,
          a_LC4_D12_aOUT, a_LC4_D12_aIN, n_6811, n_6812, n_6813, n_6814, n_6815,
          n_6816, n_6817, n_6818, a_LC8_D12_aOUT, a_LC8_D12_aIN, n_6821, n_6822,
          n_6823, n_6824, n_6825, n_6826, n_6827, a_LC6_D12_aOUT, a_LC6_D12_aIN,
          n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837,
          n_6838, a_LC7_D12_aOUT, a_LC7_D12_aIN, n_6841, n_6842, n_6843, n_6844,
          n_6845, n_6846, n_6847, n_6848, n_6849, a_N61_aCLRN, a_N61_aD, n_6856,
          n_6857, n_6858, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864,
          n_6865, n_6866, n_6867, a_N61_aCLK, a_LC2_D11_aOUT, a_LC2_D11_aIN,
          n_6871, n_6872, n_6873, n_6874, n_6875, n_6876, a_N653_aOUT, a_N653_aIN,
          n_6879, n_6880, n_6881, n_6882, n_6883, n_6884, n_6885, n_6886,
          n_6887, a_N655_aIN, n_6889, n_6890, n_6891, n_6892, n_6893, n_6894,
          n_6895, n_6896, n_6897, a_N75_aOUT, a_N75_aIN, n_6900, n_6901, n_6902,
          n_6903, n_6904, n_6905, n_6906, n_6907, a_LC3_D18_aOUT, a_LC3_D18_aIN,
          n_6910, n_6911, n_6912, n_6913, n_6914, n_6915, n_6916, a_LC2_D8_aOUT,
          a_LC2_D8_aIN, n_6919, n_6920, n_6921, n_6922, n_6923, n_6924, n_6925,
          n_6926, n_6927, n_6928, n_6929, n_6930, n_6931, n_6932, a_LC7_D8_aNOT_aOUT,
          a_LC7_D8_aNOT_aIN, n_6935, n_6936, n_6937, n_6938, n_6939, a_N656_aNOT_aOUT,
          a_N656_aNOT_aIN, n_6942, n_6943, n_6944, n_6945, n_6946, n_6947,
          n_6948, n_6949, n_6950, n_6951, a_LC5_D8_aOUT, a_LC5_D8_aIN, n_6954,
          n_6955, n_6956, n_6957, n_6958, n_6959, n_6960, n_6961, n_6962,
          n_6963, a_LC3_D12_aOUT, a_LC3_D12_aIN, n_6966, n_6967, n_6968, n_6969,
          n_6970, n_6971, n_6972, n_6973, n_6974, n_6975, a_LC5_D12_aOUT,
          a_LC5_D12_aIN, n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984,
          n_6985, n_6986, a_N63_aCLRN, a_N63_aD, n_6993, n_6994, n_6995, n_6996,
          n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, a_N63_aCLK, a_LC1_C2_aIN,
          n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011 : std_logic;

COMPONENT TRIBUF_a8251
    PORT (in1, oe  : IN std_logic; y : OUT std_logic);
END COMPONENT;

COMPONENT DFF_a8251
    PORT (d, clk, clrn, prn : IN std_logic; q : OUT std_logic);
END COMPONENT;

COMPONENT FILTER_a8251
    PORT (in1 : IN std_logic; y : OUT std_logic);
END COMPONENT;

BEGIN

PROCESS(CLK, CnD, DIN(0), DIN(1), DIN(2), DIN(3), DIN(4), DIN(5), DIN(6), DIN(7),
          EXTSYNCD, nCS, nCTS, nDSR, nRD, nRESET, nRXC, nTXC, nWR, RXD)
BEGIN
    ASSERT CLK /= 'X' OR Now = 0 ns
        REPORT "Unknown value on CLK"
        SEVERITY Warning;
    ASSERT CnD /= 'X' OR Now = 0 ns
        REPORT "Unknown value on CnD"
        SEVERITY Warning;
    ASSERT DIN(0) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(0)"
        SEVERITY Warning;
    ASSERT DIN(1) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(1)"
        SEVERITY Warning;
    ASSERT DIN(2) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(2)"
        SEVERITY Warning;
    ASSERT DIN(3) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(3)"
        SEVERITY Warning;
    ASSERT DIN(4) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(4)"
        SEVERITY Warning;
    ASSERT DIN(5) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(5)"
        SEVERITY Warning;
    ASSERT DIN(6) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(6)"
        SEVERITY Warning;
    ASSERT DIN(7) /= 'X' OR Now = 0 ns
        REPORT "Unknown value on DIN(7)"
        SEVERITY Warning;
    ASSERT EXTSYNCD /= 'X' OR Now = 0 ns
        REPORT "Unknown value on EXTSYNCD"
        SEVERITY Warning;
    ASSERT nCS /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nCS"
        SEVERITY Warning;
    ASSERT nCTS /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nCTS"
        SEVERITY Warning;
    ASSERT nDSR /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nDSR"
        SEVERITY Warning;
    ASSERT nRD /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nRD"
        SEVERITY Warning;
    ASSERT nRESET /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nRESET"
        SEVERITY Warning;
    ASSERT nRXC /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nRXC"
        SEVERITY Warning;
    ASSERT nTXC /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nTXC"
        SEVERITY Warning;
    ASSERT nWR /= 'X' OR Now = 0 ns
        REPORT "Unknown value on nWR"
        SEVERITY Warning;
    ASSERT RXD /= 'X' OR Now = 0 ns
        REPORT "Unknown value on RXD"
        SEVERITY Warning;
END PROCESS;

tribuf_2: TRIBUF_a8251
    PORT MAP (IN1 => n_83, OE => vcc, Y => DOUT(0));
tribuf_4: TRIBUF_a8251
    PORT MAP (IN1 => n_90, OE => vcc, Y => DOUT(1));
tribuf_6: TRIBUF_a8251
    PORT MAP (IN1 => n_97, OE => vcc, Y => DOUT(2));
tribuf_8: TRIBUF_a8251
    PORT MAP (IN1 => n_104, OE => vcc, Y => DOUT(3));
tribuf_10: TRIBUF_a8251
    PORT MAP (IN1 => n_111, OE => vcc, Y => DOUT(4));
tribuf_12: TRIBUF_a8251
    PORT MAP (IN1 => n_118, OE => vcc, Y => DOUT(5));
tribuf_14: TRIBUF_a8251
    PORT MAP (IN1 => n_125, OE => vcc, Y => DOUT(6));
tribuf_16: TRIBUF_a8251
    PORT MAP (IN1 => n_132, OE => vcc, Y => DOUT(7));
tribuf_18: TRIBUF_a8251
    PORT MAP (IN1 => n_139, OE => vcc, Y => TXRDY);
tribuf_20: TRIBUF_a8251
    PORT MAP (IN1 => n_146, OE => vcc, Y => TXEMPTY);
tribuf_22: TRIBUF_a8251
    PORT MAP (IN1 => n_153, OE => vcc, Y => TXD);
tribuf_24: TRIBUF_a8251
    PORT MAP (IN1 => n_160, OE => vcc, Y => SYN_BRK);
tribuf_26: TRIBUF_a8251
    PORT MAP (IN1 => n_167, OE => vcc, Y => RXRDY);
tribuf_28: TRIBUF_a8251
    PORT MAP (IN1 => n_174, OE => vcc, Y => nRTS);
tribuf_30: TRIBUF_a8251
    PORT MAP (IN1 => n_181, OE => vcc, Y => nEN);
tribuf_32: TRIBUF_a8251
    PORT MAP (IN1 => n_188, OE => vcc, Y => nDTR);
delay_33: n_83  <= TRANSPORT n_84  ;
xor2_34: n_84 <=  n_85  XOR n_89;
or1_35: n_85 <=  n_86;
and1_36: n_86 <=  n_87;
delay_37: n_87  <= TRANSPORT a_G118_aOUT  ;
and1_38: n_89 <=  gnd;
delay_39: n_90  <= TRANSPORT n_91  ;
xor2_40: n_91 <=  n_92  XOR n_96;
or1_41: n_92 <=  n_93;
and1_42: n_93 <=  n_94;
delay_43: n_94  <= TRANSPORT a_G701_aOUT  ;
and1_44: n_96 <=  gnd;
delay_45: n_97  <= TRANSPORT n_98  ;
xor2_46: n_98 <=  n_99  XOR n_103;
or1_47: n_99 <=  n_100;
and1_48: n_100 <=  n_101;
delay_49: n_101  <= TRANSPORT a_G705_aOUT  ;
and1_50: n_103 <=  gnd;
delay_51: n_104  <= TRANSPORT n_105  ;
xor2_52: n_105 <=  n_106  XOR n_110;
or1_53: n_106 <=  n_107;
and1_54: n_107 <=  n_108;
delay_55: n_108  <= TRANSPORT a_G491_aOUT  ;
and1_56: n_110 <=  gnd;
delay_57: n_111  <= TRANSPORT n_112  ;
xor2_58: n_112 <=  n_113  XOR n_117;
or1_59: n_113 <=  n_114;
and1_60: n_114 <=  n_115;
delay_61: n_115  <= TRANSPORT a_G495_aOUT  ;
and1_62: n_117 <=  gnd;
delay_63: n_118  <= TRANSPORT n_119  ;
xor2_64: n_119 <=  n_120  XOR n_124;
or1_65: n_120 <=  n_121;
and1_66: n_121 <=  n_122;
delay_67: n_122  <= TRANSPORT a_G483_aOUT  ;
and1_68: n_124 <=  gnd;
delay_69: n_125  <= TRANSPORT n_126  ;
xor2_70: n_126 <=  n_127  XOR n_131;
or1_71: n_127 <=  n_128;
and1_72: n_128 <=  n_129;
delay_73: n_129  <= TRANSPORT a_G514_aOUT  ;
and1_74: n_131 <=  gnd;
delay_75: n_132  <= TRANSPORT n_133  ;
xor2_76: n_133 <=  n_134  XOR n_138;
or1_77: n_134 <=  n_135;
and1_78: n_135 <=  n_136;
delay_79: n_136  <= TRANSPORT a_G708_aOUT  ;
and1_80: n_138 <=  gnd;
delay_81: n_139  <= TRANSPORT n_140  ;
xor2_82: n_140 <=  n_141  XOR n_145;
or1_83: n_141 <=  n_142;
and1_84: n_142 <=  n_143;
inv_85: n_143  <= TRANSPORT NOT a_STXRDY_aNOT_aQ  ;
and1_86: n_145 <=  gnd;
delay_87: n_146  <= TRANSPORT n_147  ;
xor2_88: n_147 <=  n_148  XOR n_152;
or1_89: n_148 <=  n_149;
and1_90: n_149 <=  n_150;
inv_91: n_150  <= TRANSPORT NOT a_STXEMPTY_aNOT_aQ  ;
and1_92: n_152 <=  gnd;
delay_93: n_153  <= TRANSPORT n_154  ;
xor2_94: n_154 <=  n_155  XOR n_159;
or1_95: n_155 <=  n_156;
and1_96: n_156 <=  n_157;
delay_97: n_157  <= TRANSPORT a_STXD_aOUT  ;
and1_98: n_159 <=  gnd;
delay_99: n_160  <= TRANSPORT n_161  ;
xor2_100: n_161 <=  n_162  XOR n_166;
or1_101: n_162 <=  n_163;
and1_102: n_163 <=  n_164;
delay_103: n_164  <= TRANSPORT a_SSYN_BRK_aOUT  ;
and1_104: n_166 <=  gnd;
delay_105: n_167  <= TRANSPORT n_168  ;
xor2_106: n_168 <=  n_169  XOR n_173;
or1_107: n_169 <=  n_170;
and1_108: n_170 <=  n_171;
delay_109: n_171  <= TRANSPORT a_SRXRDY_aQ  ;
and1_110: n_173 <=  gnd;
delay_111: n_174  <= TRANSPORT n_175  ;
xor2_112: n_175 <=  n_176  XOR n_180;
or1_113: n_176 <=  n_177;
and1_114: n_177 <=  n_178;
inv_115: n_178  <= TRANSPORT NOT a_SCMND_OUT_F5_G_aQ  ;
and1_116: n_180 <=  gnd;
delay_117: n_181  <= TRANSPORT n_182  ;
xor2_118: n_182 <=  n_183  XOR n_187;
or1_119: n_183 <=  n_184;
and1_120: n_184 <=  n_185;
inv_121: n_185  <= TRANSPORT NOT a_SNEN_aNOT_aOUT  ;
and1_122: n_187 <=  gnd;
delay_123: n_188  <= TRANSPORT n_189  ;
xor2_124: n_189 <=  n_190  XOR n_194;
or1_125: n_190 <=  n_191;
and1_126: n_191 <=  n_192;
inv_127: n_192  <= TRANSPORT NOT a_SCMND_OUT_F1_G_aQ  ;
and1_128: n_194 <=  gnd;
delay_129: a_N580_aNOT_aOUT  <= TRANSPORT a_N580_aNOT_aIN  ;
xor2_130: a_N580_aNOT_aIN <=  n_197  XOR n_203;
or1_131: n_197 <=  n_198;
and2_132: n_198 <=  n_199  AND n_201;
delay_133: n_199  <= TRANSPORT a_N607_aOUT  ;
delay_134: n_201  <= TRANSPORT a_LC1_C2_aOUT  ;
and1_135: n_203 <=  gnd;
dff_136: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F3_G_aD, CLK => a_SMODE_OUT_F3_G_aCLK, CLRN => a_SMODE_OUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F3_G_aQ);
delay_137: a_SMODE_OUT_F3_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_138: a_SMODE_OUT_F3_G_aD <=  n_212  XOR n_221;
or2_139: n_212 <=  n_213  OR n_215;
and1_140: n_213 <=  n_214;
delay_141: n_214  <= TRANSPORT a_N580_aNOT_aOUT  ;
and3_142: n_215 <=  n_216  AND n_218  AND n_220;
delay_143: n_216  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_144: n_218  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_145: n_220  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_146: n_221 <=  gnd;
delay_147: n_222  <= TRANSPORT CLK  ;
filter_148: FILTER_a8251
    PORT MAP (IN1 => n_222, Y => a_SMODE_OUT_F3_G_aCLK);
delay_149: a_LC2_C16_aOUT  <= TRANSPORT a_LC2_C16_aIN  ;
xor2_150: a_LC2_C16_aIN <=  n_227  XOR n_234;
or1_151: n_227 <=  n_228;
and3_152: n_228 <=  n_229  AND n_231  AND n_233;
delay_153: n_229  <= TRANSPORT a_N1189_aOUT  ;
delay_154: n_231  <= TRANSPORT DIN(2)  ;
delay_155: n_233  <= TRANSPORT a_LC1_C2_aOUT  ;
and1_156: n_234 <=  gnd;
dff_157: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F2_G_aD, CLK => a_SMODE_OUT_F2_G_aCLK, CLRN => a_SMODE_OUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F2_G_aQ);
delay_158: a_SMODE_OUT_F2_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_159: a_SMODE_OUT_F2_G_aD <=  n_242  XOR n_250;
or2_160: n_242 <=  n_243  OR n_246;
and2_161: n_243 <=  n_244  AND n_245;
delay_162: n_244  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_163: n_245  <= TRANSPORT a_LC2_C16_aOUT  ;
and3_164: n_246 <=  n_247  AND n_248  AND n_249;
delay_165: n_247  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_166: n_248  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_167: n_249  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_168: n_250 <=  gnd;
delay_169: n_251  <= TRANSPORT CLK  ;
filter_170: FILTER_a8251
    PORT MAP (IN1 => n_251, Y => a_SMODE_OUT_F2_G_aCLK);
dff_171: DFF_a8251
    PORT MAP ( D => a_N1804_aD, CLK => a_N1804_aCLK, CLRN => a_N1804_aCLRN,
          PRN => vcc, Q => a_N1804_aQ);
delay_172: a_N1804_aCLRN  <= TRANSPORT nRESET  ;
xor2_173: a_N1804_aD <=  n_260  XOR n_264;
or1_174: n_260 <=  n_261;
and1_175: n_261 <=  n_262;
delay_176: n_262  <= TRANSPORT a_N1807_aQ  ;
and1_177: n_264 <=  gnd;
delay_178: n_265  <= TRANSPORT CLK  ;
filter_179: FILTER_a8251
    PORT MAP (IN1 => n_265, Y => a_N1804_aCLK);
dff_180: DFF_a8251
    PORT MAP ( D => a_N1807_aD, CLK => a_N1807_aCLK, CLRN => a_N1807_aCLRN,
          PRN => vcc, Q => a_N1807_aQ);
delay_181: a_N1807_aCLRN  <= TRANSPORT nRESET  ;
xor2_182: a_N1807_aD <=  n_273  XOR n_281;
or1_183: n_273 <=  n_274;
and3_184: n_274 <=  n_275  AND n_277  AND n_279;
inv_185: n_275  <= TRANSPORT NOT nWR  ;
delay_186: n_277  <= TRANSPORT CnD  ;
inv_187: n_279  <= TRANSPORT NOT nCS  ;
and1_188: n_281 <=  gnd;
delay_189: n_282  <= TRANSPORT CLK  ;
filter_190: FILTER_a8251
    PORT MAP (IN1 => n_282, Y => a_N1807_aCLK);
delay_191: a_LC8_C7_aOUT  <= TRANSPORT a_LC8_C7_aIN  ;
xor2_192: a_LC8_C7_aIN <=  n_286  XOR n_299;
or2_193: n_286 <=  n_287  OR n_294;
and3_194: n_287 <=  n_288  AND n_290  AND n_292;
inv_195: n_288  <= TRANSPORT NOT a_LC1_C7_aNOT_aOUT  ;
inv_196: n_290  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_197: n_292  <= TRANSPORT a_SCMND_OUT_F4_G_aQ  ;
and3_198: n_294 <=  n_295  AND n_297  AND n_298;
delay_199: n_295  <= TRANSPORT DIN(4)  ;
delay_200: n_297  <= TRANSPORT a_LC1_C7_aNOT_aOUT  ;
inv_201: n_298  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
and1_202: n_299 <=  gnd;
dff_203: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F4_G_aD, CLK => a_SCMND_OUT_F4_G_aCLK, CLRN => a_SCMND_OUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F4_G_aQ);
delay_204: a_SCMND_OUT_F4_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_205: a_SCMND_OUT_F4_G_aD <=  n_306  XOR n_310;
or1_206: n_306 <=  n_307;
and2_207: n_307 <=  n_308  AND n_309;
delay_208: n_308  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_209: n_309  <= TRANSPORT a_LC8_C7_aOUT  ;
and1_210: n_310 <=  gnd;
delay_211: n_311  <= TRANSPORT CLK  ;
filter_212: FILTER_a8251
    PORT MAP (IN1 => n_311, Y => a_SCMND_OUT_F4_G_aCLK);
delay_213: a_N101_aOUT  <= TRANSPORT a_N101_aIN  ;
xor2_214: a_N101_aIN <=  n_315  XOR n_321;
or1_215: n_315 <=  n_316;
and2_216: n_316 <=  n_317  AND n_319;
delay_217: n_317  <= TRANSPORT a_N1757_aQ  ;
inv_218: n_319  <= TRANSPORT NOT a_N1756_aQ  ;
and1_219: n_321 <=  gnd;
delay_220: a_N227_aNOT_aOUT  <= TRANSPORT a_N227_aNOT_aIN  ;
xor2_221: a_N227_aNOT_aIN <=  n_324  XOR n_333;
or1_222: n_324 <=  n_325;
and4_223: n_325 <=  n_326  AND n_328  AND n_330  AND n_331;
delay_224: n_326  <= TRANSPORT a_N130_aNOT_aOUT  ;
delay_225: n_328  <= TRANSPORT a_N1165_aOUT  ;
delay_226: n_330  <= TRANSPORT a_N101_aOUT  ;
inv_227: n_331  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_228: n_333 <=  gnd;
delay_229: a_LC5_C20_aOUT  <= TRANSPORT a_LC5_C20_aIN  ;
xor2_230: a_LC5_C20_aIN <=  n_336  XOR n_346;
or2_231: n_336 <=  n_337  OR n_342;
and3_232: n_337 <=  n_338  AND n_340  AND n_341;
delay_233: n_338  <= TRANSPORT a_N1754_aQ  ;
inv_234: n_340  <= TRANSPORT NOT a_N1757_aQ  ;
inv_235: n_341  <= TRANSPORT NOT a_N1756_aQ  ;
and3_236: n_342 <=  n_343  AND n_344  AND n_345;
inv_237: n_343  <= TRANSPORT NOT a_N227_aNOT_aOUT  ;
delay_238: n_344  <= TRANSPORT a_N1757_aQ  ;
inv_239: n_345  <= TRANSPORT NOT a_N1756_aQ  ;
and1_240: n_346 <=  gnd;
delay_241: a_N239_aOUT  <= TRANSPORT a_N239_aIN  ;
xor2_242: a_N239_aIN <=  n_349  XOR n_359;
or2_243: n_349 <=  n_350  OR n_354;
and3_244: n_350 <=  n_351  AND n_352  AND n_353;
delay_245: n_351  <= TRANSPORT a_N1165_aOUT  ;
delay_246: n_352  <= TRANSPORT a_N1757_aQ  ;
delay_247: n_353  <= TRANSPORT a_N1756_aQ  ;
and3_248: n_354 <=  n_355  AND n_356  AND n_358;
delay_249: n_355  <= TRANSPORT a_N1165_aOUT  ;
delay_250: n_356  <= TRANSPORT a_SMODE_OUT_F7_G_aQ  ;
delay_251: n_358  <= TRANSPORT a_N1756_aQ  ;
and1_252: n_359 <=  gnd;
dff_253: DFF_a8251
    PORT MAP ( D => a_N1754_aD, CLK => a_N1754_aCLK, CLRN => a_N1754_aCLRN,
          PRN => vcc, Q => a_N1754_aQ);
delay_254: a_N1754_aCLRN  <= TRANSPORT nRESET  ;
xor2_255: a_N1754_aD <=  n_366  XOR n_373;
or2_256: n_366 <=  n_367  OR n_370;
and2_257: n_367 <=  n_368  AND n_369;
delay_258: n_368  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_259: n_369  <= TRANSPORT a_LC5_C20_aOUT  ;
and2_260: n_370 <=  n_371  AND n_372;
delay_261: n_371  <= TRANSPORT a_N1189_aOUT  ;
delay_262: n_372  <= TRANSPORT a_N239_aOUT  ;
and1_263: n_373 <=  gnd;
delay_264: n_374  <= TRANSPORT CLK  ;
filter_265: FILTER_a8251
    PORT MAP (IN1 => n_374, Y => a_N1754_aCLK);
delay_266: a_N236_aOUT  <= TRANSPORT a_N236_aIN  ;
xor2_267: a_N236_aIN <=  n_378  XOR n_388;
or2_268: n_378 <=  n_379  OR n_384;
and4_269: n_379 <=  n_380  AND n_381  AND n_382  AND n_383;
delay_270: n_380  <= TRANSPORT a_N1189_aOUT  ;
inv_271: n_381  <= TRANSPORT NOT a_SMODE_OUT_F7_G_aQ  ;
inv_272: n_382  <= TRANSPORT NOT a_N1757_aQ  ;
delay_273: n_383  <= TRANSPORT a_N1756_aQ  ;
and3_274: n_384 <=  n_385  AND n_386  AND n_387;
inv_275: n_385  <= TRANSPORT NOT a_N1189_aOUT  ;
delay_276: n_386  <= TRANSPORT a_N1757_aQ  ;
delay_277: n_387  <= TRANSPORT a_N1756_aQ  ;
and1_278: n_388 <=  gnd;
dff_279: DFF_a8251
    PORT MAP ( D => a_N1757_aD, CLK => a_N1757_aCLK, CLRN => a_N1757_aCLRN,
          PRN => vcc, Q => a_N1757_aQ);
delay_280: a_N1757_aCLRN  <= TRANSPORT nRESET  ;
xor2_281: a_N1757_aD <=  n_395  XOR n_401;
or2_282: n_395 <=  n_396  OR n_399;
and2_283: n_396 <=  n_397  AND n_398;
delay_284: n_397  <= TRANSPORT a_N1165_aOUT  ;
delay_285: n_398  <= TRANSPORT a_N236_aOUT  ;
and1_286: n_399 <=  n_400;
inv_287: n_400  <= TRANSPORT NOT a_N1034_aNOT_aOUT  ;
and1_288: n_401 <=  gnd;
delay_289: n_402  <= TRANSPORT CLK  ;
filter_290: FILTER_a8251
    PORT MAP (IN1 => n_402, Y => a_N1757_aCLK);
delay_291: a_N235_aNOT_aOUT  <= TRANSPORT a_N235_aNOT_aIN  ;
xor2_292: a_N235_aNOT_aIN <=  n_406  XOR n_412;
or1_293: n_406 <=  n_407;
and4_294: n_407 <=  n_408  AND n_409  AND n_410  AND n_411;
inv_295: n_408  <= TRANSPORT NOT a_N1189_aOUT  ;
delay_296: n_409  <= TRANSPORT a_N1165_aOUT  ;
inv_297: n_410  <= TRANSPORT NOT a_N1757_aQ  ;
delay_298: n_411  <= TRANSPORT a_N1756_aQ  ;
and1_299: n_412 <=  gnd;
dff_300: DFF_a8251
    PORT MAP ( D => a_N1756_aD, CLK => a_N1756_aCLK, CLRN => a_N1756_aCLRN,
          PRN => vcc, Q => a_N1756_aQ);
delay_301: a_N1756_aCLRN  <= TRANSPORT nRESET  ;
xor2_302: a_N1756_aD <=  n_419  XOR n_427;
or3_303: n_419 <=  n_420  OR n_423  OR n_425;
and2_304: n_420 <=  n_421  AND n_422;
delay_305: n_421  <= TRANSPORT a_N1165_aOUT  ;
delay_306: n_422  <= TRANSPORT a_N236_aOUT  ;
and1_307: n_423 <=  n_424;
delay_308: n_424  <= TRANSPORT a_N235_aNOT_aOUT  ;
and1_309: n_425 <=  n_426;
delay_310: n_426  <= TRANSPORT a_N227_aNOT_aOUT  ;
and1_311: n_427 <=  gnd;
delay_312: n_428  <= TRANSPORT CLK  ;
filter_313: FILTER_a8251
    PORT MAP (IN1 => n_428, Y => a_N1756_aCLK);
dff_314: DFF_a8251
    PORT MAP ( D => a_N1806_aD, CLK => a_N1806_aCLK, CLRN => a_N1806_aCLRN,
          PRN => vcc, Q => a_N1806_aQ);
delay_315: a_N1806_aCLRN  <= TRANSPORT nRESET  ;
xor2_316: a_N1806_aD <=  n_437  XOR n_441;
or1_317: n_437 <=  n_438;
and1_318: n_438 <=  n_439;
delay_319: n_439  <= TRANSPORT a_N1808_aQ  ;
and1_320: n_441 <=  gnd;
delay_321: n_442  <= TRANSPORT CLK  ;
filter_322: FILTER_a8251
    PORT MAP (IN1 => n_442, Y => a_N1806_aCLK);
dff_323: DFF_a8251
    PORT MAP ( D => a_N1808_aD, CLK => a_N1808_aCLK, CLRN => a_N1808_aCLRN,
          PRN => vcc, Q => a_N1808_aQ);
delay_324: a_N1808_aCLRN  <= TRANSPORT nRESET  ;
xor2_325: a_N1808_aD <=  n_450  XOR n_457;
or1_326: n_450 <=  n_451;
and4_327: n_451 <=  n_452  AND n_454  AND n_455  AND n_456;
delay_328: n_452  <= TRANSPORT mode_cmplt_aOUT  ;
inv_329: n_454  <= TRANSPORT NOT nWR  ;
delay_330: n_455  <= TRANSPORT CnD  ;
inv_331: n_456  <= TRANSPORT NOT nCS  ;
and1_332: n_457 <=  gnd;
delay_333: n_458  <= TRANSPORT CLK  ;
filter_334: FILTER_a8251
    PORT MAP (IN1 => n_458, Y => a_N1808_aCLK);
dff_335: DFF_a8251
    PORT MAP ( D => a_N1898_aD, CLK => a_N1898_aCLK, CLRN => a_N1898_aCLRN,
          PRN => vcc, Q => a_N1898_aQ);
delay_336: a_N1898_aCLRN  <= TRANSPORT nRESET  ;
xor2_337: a_N1898_aD <=  n_468  XOR n_471;
or1_338: n_468 <=  n_469;
and1_339: n_469 <=  n_470;
delay_340: n_470  <= TRANSPORT a_SCMND_OUT_F4_G_aQ  ;
and1_341: n_471 <=  gnd;
delay_342: n_472  <= TRANSPORT nRXC  ;
filter_343: FILTER_a8251
    PORT MAP (IN1 => n_472, Y => a_N1898_aCLK);
dff_344: DFF_a8251
    PORT MAP ( D => a_N1897_aD, CLK => a_N1897_aCLK, CLRN => a_N1897_aCLRN,
          PRN => vcc, Q => a_N1897_aQ);
delay_345: a_N1897_aCLRN  <= TRANSPORT nRESET  ;
xor2_346: a_N1897_aD <=  n_482  XOR n_485;
or1_347: n_482 <=  n_483;
and1_348: n_483 <=  n_484;
delay_349: n_484  <= TRANSPORT a_N1898_aQ  ;
and1_350: n_485 <=  gnd;
delay_351: n_486  <= TRANSPORT nRXC  ;
filter_352: FILTER_a8251
    PORT MAP (IN1 => n_486, Y => a_N1897_aCLK);
delay_353: a_N310_aNOT_aOUT  <= TRANSPORT a_N310_aNOT_aIN  ;
xor2_354: a_N310_aNOT_aIN <=  n_490  XOR n_500;
or2_355: n_490 <=  n_491  OR n_496;
and2_356: n_491 <=  n_492  AND n_494;
inv_357: n_492  <= TRANSPORT NOT a_N296_aNOT_aOUT  ;
delay_358: n_494  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and2_359: n_496 <=  n_497  AND n_498;
inv_360: n_497  <= TRANSPORT NOT a_N296_aNOT_aOUT  ;
delay_361: n_498  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and1_362: n_500 <=  gnd;
delay_363: a_LC3_B16_aOUT  <= TRANSPORT a_LC3_B16_aIN  ;
xor2_364: a_LC3_B16_aIN <=  n_503  XOR n_516;
or2_365: n_503 <=  n_504  OR n_511;
and3_366: n_504 <=  n_505  AND n_507  AND n_509;
delay_367: n_505  <= TRANSPORT a_N1107_aOUT  ;
delay_368: n_507  <= TRANSPORT a_N414_aQ  ;
inv_369: n_509  <= TRANSPORT NOT a_N413_aQ  ;
and3_370: n_511 <=  n_512  AND n_514  AND n_515;
delay_371: n_512  <= TRANSPORT a_N298_aOUT  ;
inv_372: n_514  <= TRANSPORT NOT a_N414_aQ  ;
inv_373: n_515  <= TRANSPORT NOT a_N413_aQ  ;
and1_374: n_516 <=  gnd;
dff_375: DFF_a8251
    PORT MAP ( D => a_N411_aD, CLK => a_N411_aCLK, CLRN => a_N411_aCLRN, PRN => vcc,
          Q => a_N411_aQ);
delay_376: a_N411_aCLRN  <= TRANSPORT nRESET  ;
xor2_377: a_N411_aD <=  n_524  XOR n_533;
or2_378: n_524 <=  n_525  OR n_529;
and2_379: n_525 <=  n_526  AND n_528;
delay_380: n_526  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_381: n_528  <= TRANSPORT a_N310_aNOT_aOUT  ;
and3_382: n_529 <=  n_530  AND n_531  AND n_532;
delay_383: n_530  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_384: n_531  <= TRANSPORT a_LC3_B16_aOUT  ;
delay_385: n_532  <= TRANSPORT a_N411_aQ  ;
and1_386: n_533 <=  gnd;
inv_387: n_534  <= TRANSPORT NOT nTXC  ;
filter_388: FILTER_a8251
    PORT MAP (IN1 => n_534, Y => a_N411_aCLK);
delay_389: a_LC5_B18_aOUT  <= TRANSPORT a_LC5_B18_aIN  ;
xor2_390: a_LC5_B18_aIN <=  n_539  XOR n_550;
or2_391: n_539 <=  n_540  OR n_545;
and2_392: n_540 <=  n_541  AND n_543;
delay_393: n_541  <= TRANSPORT a_N470_aOUT  ;
delay_394: n_543  <= TRANSPORT a_N869_aQ  ;
and2_395: n_545 <=  n_546  AND n_548;
delay_396: n_546  <= TRANSPORT a_LC2_B11_aOUT  ;
delay_397: n_548  <= TRANSPORT a_N606_aQ  ;
and1_398: n_550 <=  gnd;
delay_399: a_N179_aOUT  <= TRANSPORT a_N179_aIN  ;
xor2_400: a_N179_aIN <=  n_553  XOR n_563;
or2_401: n_553 <=  n_554  OR n_559;
and2_402: n_554 <=  n_555  AND n_557;
delay_403: n_555  <= TRANSPORT a_SSYNC2_F0_G_aQ  ;
delay_404: n_557  <= TRANSPORT a_N729_aQ  ;
and2_405: n_559 <=  n_560  AND n_561;
inv_406: n_560  <= TRANSPORT NOT a_N729_aQ  ;
delay_407: n_561  <= TRANSPORT a_SSYNC1_F0_G_aQ  ;
and1_408: n_563 <=  gnd;
delay_409: a_N1093_aNOT_aOUT  <= TRANSPORT a_N1093_aNOT_aIN  ;
xor2_410: a_N1093_aNOT_aIN <=  n_566  XOR n_575;
or2_411: n_566 <=  n_567  OR n_571;
and2_412: n_567 <=  n_568  AND n_570;
inv_413: n_568  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_414: n_570  <= TRANSPORT a_N179_aOUT  ;
and2_415: n_571 <=  n_572  AND n_573;
delay_416: n_572  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_417: n_573  <= TRANSPORT a_N2031_aQ  ;
and1_418: n_575 <=  gnd;
dff_419: DFF_a8251
    PORT MAP ( D => a_N869_aD, CLK => a_N869_aCLK, CLRN => a_N869_aCLRN, PRN => vcc,
          Q => a_N869_aQ);
delay_420: a_N869_aCLRN  <= TRANSPORT nRESET  ;
xor2_421: a_N869_aD <=  n_582  XOR n_592;
or2_422: n_582 <=  n_583  OR n_588;
and3_423: n_583 <=  n_584  AND n_585  AND n_587;
delay_424: n_584  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_425: n_585  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_426: n_587  <= TRANSPORT a_LC5_B18_aOUT  ;
and3_427: n_588 <=  n_589  AND n_590  AND n_591;
delay_428: n_589  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_429: n_590  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_430: n_591  <= TRANSPORT a_N1093_aNOT_aOUT  ;
and1_431: n_592 <=  gnd;
inv_432: n_593  <= TRANSPORT NOT nTXC  ;
filter_433: FILTER_a8251
    PORT MAP (IN1 => n_593, Y => a_N869_aCLK);
dff_434: DFF_a8251
    PORT MAP ( D => a_N1904_aD, CLK => a_N1904_aCLK, CLRN => a_N1904_aCLRN,
          PRN => vcc, Q => a_N1904_aQ);
delay_435: a_N1904_aCLRN  <= TRANSPORT nRESET  ;
xor2_436: a_N1904_aD <=  n_603  XOR n_609;
or1_437: n_603 <=  n_604;
and4_438: n_604 <=  n_605  AND n_606  AND n_607  AND n_608;
delay_439: n_605  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_440: n_606  <= TRANSPORT a_N1754_aQ  ;
inv_441: n_607  <= TRANSPORT NOT a_N1757_aQ  ;
inv_442: n_608  <= TRANSPORT NOT a_N1756_aQ  ;
and1_443: n_609 <=  gnd;
delay_444: n_610  <= TRANSPORT nTXC  ;
filter_445: FILTER_a8251
    PORT MAP (IN1 => n_610, Y => a_N1904_aCLK);
dff_446: DFF_a8251
    PORT MAP ( D => a_N1903_aD, CLK => a_N1903_aCLK, CLRN => a_N1903_aCLRN,
          PRN => vcc, Q => a_N1903_aQ);
delay_447: a_N1903_aCLRN  <= TRANSPORT nRESET  ;
xor2_448: a_N1903_aD <=  n_619  XOR n_622;
or1_449: n_619 <=  n_620;
and1_450: n_620 <=  n_621;
delay_451: n_621  <= TRANSPORT a_N1904_aQ  ;
and1_452: n_622 <=  gnd;
delay_453: n_623  <= TRANSPORT nTXC  ;
filter_454: FILTER_a8251
    PORT MAP (IN1 => n_623, Y => a_N1903_aCLK);
delay_455: a_LC6_C3_aOUT  <= TRANSPORT a_LC6_C3_aIN  ;
xor2_456: a_LC6_C3_aIN <=  n_627  XOR n_633;
or1_457: n_627 <=  n_628;
and3_458: n_628 <=  n_629  AND n_630  AND n_632;
delay_459: n_629  <= TRANSPORT a_N1189_aOUT  ;
inv_460: n_630  <= TRANSPORT NOT a_N1123_aNOT_aOUT  ;
delay_461: n_632  <= TRANSPORT DIN(4)  ;
and1_462: n_633 <=  gnd;
dff_463: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F4_G_aD, CLK => a_SMODE_OUT_F4_G_aCLK, CLRN => a_SMODE_OUT_F4_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F4_G_aQ);
delay_464: a_SMODE_OUT_F4_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_465: a_SMODE_OUT_F4_G_aD <=  n_641  XOR n_649;
or2_466: n_641 <=  n_642  OR n_646;
and3_467: n_642 <=  n_643  AND n_644  AND n_645;
delay_468: n_643  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_469: n_644  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_470: n_645  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_471: n_646 <=  n_647  AND n_648;
delay_472: n_647  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_473: n_648  <= TRANSPORT a_LC6_C3_aOUT  ;
and1_474: n_649 <=  gnd;
delay_475: n_650  <= TRANSPORT CLK  ;
filter_476: FILTER_a8251
    PORT MAP (IN1 => n_650, Y => a_SMODE_OUT_F4_G_aCLK);
delay_477: a_LC1_C3_aOUT  <= TRANSPORT a_LC1_C3_aIN  ;
xor2_478: a_LC1_C3_aIN <=  n_654  XOR n_661;
or1_479: n_654 <=  n_655;
and4_480: n_655 <=  n_656  AND n_657  AND n_658  AND n_659;
delay_481: n_656  <= TRANSPORT a_N1189_aOUT  ;
delay_482: n_657  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_483: n_658  <= TRANSPORT NOT a_N1123_aNOT_aOUT  ;
delay_484: n_659  <= TRANSPORT DIN(6)  ;
and1_485: n_661 <=  gnd;
dff_486: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F6_G_aD, CLK => a_SMODE_OUT_F6_G_aCLK, CLRN => a_SMODE_OUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F6_G_aQ);
delay_487: a_SMODE_OUT_F6_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_488: a_SMODE_OUT_F6_G_aD <=  n_668  XOR n_676;
or2_489: n_668 <=  n_669  OR n_672;
and2_490: n_669 <=  n_670  AND n_671;
delay_491: n_670  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_492: n_671  <= TRANSPORT a_LC1_C3_aOUT  ;
and3_493: n_672 <=  n_673  AND n_674  AND n_675;
delay_494: n_673  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_495: n_674  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_496: n_675  <= TRANSPORT a_SMODE_OUT_F6_G_aQ  ;
and1_497: n_676 <=  gnd;
delay_498: n_677  <= TRANSPORT CLK  ;
filter_499: FILTER_a8251
    PORT MAP (IN1 => n_677, Y => a_SMODE_OUT_F6_G_aCLK);
dff_500: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F6_G_aD, CLK => a_SCMND_OUT_F6_G_aCLK, CLRN => a_SCMND_OUT_F6_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F6_G_aQ);
delay_501: a_SCMND_OUT_F6_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_502: a_SCMND_OUT_F6_G_aD <=  n_686  XOR n_696;
or2_503: n_686 <=  n_687  OR n_692;
and3_504: n_687 <=  n_688  AND n_689  AND n_691;
delay_505: n_688  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_506: n_689  <= TRANSPORT NOT a_N701_aNOT_aOUT  ;
delay_507: n_691  <= TRANSPORT a_SCMND_OUT_F6_G_aQ  ;
and3_508: n_692 <=  n_693  AND n_694  AND n_695;
delay_509: n_693  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_510: n_694  <= TRANSPORT a_N701_aNOT_aOUT  ;
delay_511: n_695  <= TRANSPORT DIN(6)  ;
and1_512: n_696 <=  gnd;
delay_513: n_697  <= TRANSPORT CLK  ;
filter_514: FILTER_a8251
    PORT MAP (IN1 => n_697, Y => a_SCMND_OUT_F6_G_aCLK);
dff_515: DFF_a8251
    PORT MAP ( D => a_N1895_aD, CLK => a_N1895_aCLK, CLRN => a_N1895_aCLRN,
          PRN => vcc, Q => a_N1895_aQ);
delay_516: a_N1895_aCLRN  <= TRANSPORT nRESET  ;
xor2_517: a_N1895_aD <=  n_706  XOR n_709;
or1_518: n_706 <=  n_707;
and1_519: n_707 <=  n_708;
delay_520: n_708  <= TRANSPORT a_SCMND_OUT_F6_G_aQ  ;
and1_521: n_709 <=  gnd;
delay_522: n_710  <= TRANSPORT CLK  ;
filter_523: FILTER_a8251
    PORT MAP (IN1 => n_710, Y => a_N1895_aCLK);
dff_524: DFF_a8251
    PORT MAP ( D => a_N1811_aD, CLK => a_N1811_aCLK, CLRN => a_N1811_aCLRN,
          PRN => vcc, Q => a_N1811_aQ);
delay_525: a_N1811_aCLRN  <= TRANSPORT nRESET  ;
xor2_526: a_N1811_aD <=  n_719  XOR n_723;
or1_527: n_719 <=  n_720;
and1_528: n_720 <=  n_721;
delay_529: n_721  <= TRANSPORT a_N1812_aQ  ;
and1_530: n_723 <=  gnd;
delay_531: n_724  <= TRANSPORT nTXC  ;
filter_532: FILTER_a8251
    PORT MAP (IN1 => n_724, Y => a_N1811_aCLK);
delay_533: a_N100_aOUT  <= TRANSPORT a_N100_aIN  ;
xor2_534: a_N100_aIN <=  n_728  XOR n_734;
or1_535: n_728 <=  n_729;
and3_536: n_729 <=  n_730  AND n_732  AND n_733;
inv_537: n_730  <= TRANSPORT NOT a_LC5_C13_aOUT  ;
inv_538: n_732  <= TRANSPORT NOT CnD  ;
delay_539: n_733  <= TRANSPORT nRESET  ;
and1_540: n_734 <=  gnd;
dff_541: DFF_a8251
    PORT MAP ( D => a_N1812_aD, CLK => a_N1812_aCLK, CLRN => a_N1812_aCLRN,
          PRN => vcc, Q => a_N1812_aQ);
delay_542: a_N1812_aCLRN  <= TRANSPORT nRESET  ;
xor2_543: a_N1812_aD <=  n_741  XOR n_748;
or1_544: n_741 <=  n_742;
and4_545: n_742 <=  n_743  AND n_744  AND n_745  AND n_747;
inv_546: n_743  <= TRANSPORT NOT nWR  ;
delay_547: n_744  <= TRANSPORT a_N100_aOUT  ;
delay_548: n_745  <= TRANSPORT nRD  ;
inv_549: n_747  <= TRANSPORT NOT nCS  ;
and1_550: n_748 <=  gnd;
delay_551: n_749  <= TRANSPORT nTXC  ;
filter_552: FILTER_a8251
    PORT MAP (IN1 => n_749, Y => a_N1812_aCLK);
delay_553: a_LC8_B20_aOUT  <= TRANSPORT a_LC8_B20_aIN  ;
xor2_554: a_LC8_B20_aIN <=  n_753  XOR n_771;
or4_555: n_753 <=  n_754  OR n_759  OR n_763  OR n_767;
and3_556: n_754 <=  n_755  AND n_756  AND n_757;
delay_557: n_755  <= TRANSPORT a_N1114_aNOT_aOUT  ;
inv_558: n_756  <= TRANSPORT NOT a_N2031_aQ  ;
inv_559: n_757  <= TRANSPORT NOT a_SMODE_OUT_F5_G_aQ  ;
and3_560: n_759 <=  n_760  AND n_761  AND n_762;
delay_561: n_760  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_562: n_761  <= TRANSPORT a_N2031_aQ  ;
delay_563: n_762  <= TRANSPORT a_SMODE_OUT_F5_G_aQ  ;
and3_564: n_763 <=  n_764  AND n_765  AND n_766;
inv_565: n_764  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_566: n_765  <= TRANSPORT a_SMODE_OUT_F5_G_aQ  ;
delay_567: n_766  <= TRANSPORT a_N179_aOUT  ;
and3_568: n_767 <=  n_768  AND n_769  AND n_770;
inv_569: n_768  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
inv_570: n_769  <= TRANSPORT NOT a_SMODE_OUT_F5_G_aQ  ;
inv_571: n_770  <= TRANSPORT NOT a_N179_aOUT  ;
and1_572: n_771 <=  gnd;
delay_573: a_LC4_B2_aOUT  <= TRANSPORT a_LC4_B2_aIN  ;
xor2_574: a_LC4_B2_aIN <=  n_774  XOR n_819;
or8_575: n_774 <=  n_775  OR n_784  OR n_789  OR n_794  OR n_799  OR n_804
           OR n_809  OR n_814;
and4_576: n_775 <=  n_776  AND n_778  AND n_780  AND n_782;
delay_577: n_776  <= TRANSPORT a_N1108_aNOT_aOUT  ;
inv_578: n_778  <= TRANSPORT NOT a_N1099_aNOT_aOUT  ;
delay_579: n_780  <= TRANSPORT a_N1098_aNOT_aOUT  ;
delay_580: n_782  <= TRANSPORT a_N1097_aNOT_aOUT  ;
and4_581: n_784 <=  n_785  AND n_786  AND n_787  AND n_788;
inv_582: n_785  <= TRANSPORT NOT a_N1108_aNOT_aOUT  ;
delay_583: n_786  <= TRANSPORT a_N1099_aNOT_aOUT  ;
delay_584: n_787  <= TRANSPORT a_N1098_aNOT_aOUT  ;
delay_585: n_788  <= TRANSPORT a_N1097_aNOT_aOUT  ;
and4_586: n_789 <=  n_790  AND n_791  AND n_792  AND n_793;
inv_587: n_790  <= TRANSPORT NOT a_N1108_aNOT_aOUT  ;
inv_588: n_791  <= TRANSPORT NOT a_N1099_aNOT_aOUT  ;
inv_589: n_792  <= TRANSPORT NOT a_N1098_aNOT_aOUT  ;
delay_590: n_793  <= TRANSPORT a_N1097_aNOT_aOUT  ;
and4_591: n_794 <=  n_795  AND n_796  AND n_797  AND n_798;
delay_592: n_795  <= TRANSPORT a_N1108_aNOT_aOUT  ;
delay_593: n_796  <= TRANSPORT a_N1099_aNOT_aOUT  ;
inv_594: n_797  <= TRANSPORT NOT a_N1098_aNOT_aOUT  ;
delay_595: n_798  <= TRANSPORT a_N1097_aNOT_aOUT  ;
and4_596: n_799 <=  n_800  AND n_801  AND n_802  AND n_803;
delay_597: n_800  <= TRANSPORT a_N1108_aNOT_aOUT  ;
inv_598: n_801  <= TRANSPORT NOT a_N1099_aNOT_aOUT  ;
inv_599: n_802  <= TRANSPORT NOT a_N1098_aNOT_aOUT  ;
inv_600: n_803  <= TRANSPORT NOT a_N1097_aNOT_aOUT  ;
and4_601: n_804 <=  n_805  AND n_806  AND n_807  AND n_808;
inv_602: n_805  <= TRANSPORT NOT a_N1108_aNOT_aOUT  ;
delay_603: n_806  <= TRANSPORT a_N1099_aNOT_aOUT  ;
inv_604: n_807  <= TRANSPORT NOT a_N1098_aNOT_aOUT  ;
inv_605: n_808  <= TRANSPORT NOT a_N1097_aNOT_aOUT  ;
and4_606: n_809 <=  n_810  AND n_811  AND n_812  AND n_813;
inv_607: n_810  <= TRANSPORT NOT a_N1108_aNOT_aOUT  ;
inv_608: n_811  <= TRANSPORT NOT a_N1099_aNOT_aOUT  ;
delay_609: n_812  <= TRANSPORT a_N1098_aNOT_aOUT  ;
inv_610: n_813  <= TRANSPORT NOT a_N1097_aNOT_aOUT  ;
and4_611: n_814 <=  n_815  AND n_816  AND n_817  AND n_818;
delay_612: n_815  <= TRANSPORT a_N1108_aNOT_aOUT  ;
delay_613: n_816  <= TRANSPORT a_N1099_aNOT_aOUT  ;
delay_614: n_817  <= TRANSPORT a_N1098_aNOT_aOUT  ;
inv_615: n_818  <= TRANSPORT NOT a_N1097_aNOT_aOUT  ;
and1_616: n_819 <=  gnd;
delay_617: a_LC7_B2_aOUT  <= TRANSPORT a_LC7_B2_aIN  ;
xor2_618: a_LC7_B2_aIN <=  n_822  XOR n_866;
or8_619: n_822 <=  n_823  OR n_831  OR n_836  OR n_841  OR n_846  OR n_851
           OR n_856  OR n_861;
and4_620: n_823 <=  n_824  AND n_826  AND n_828  AND n_830;
delay_621: n_824  <= TRANSPORT a_N1096_aNOT_aOUT  ;
delay_622: n_826  <= TRANSPORT a_N1095_aNOT_aOUT  ;
delay_623: n_828  <= TRANSPORT a_N1094_aNOT_aOUT  ;
delay_624: n_830  <= TRANSPORT a_LC4_B2_aOUT  ;
and4_625: n_831 <=  n_832  AND n_833  AND n_834  AND n_835;
inv_626: n_832  <= TRANSPORT NOT a_N1096_aNOT_aOUT  ;
inv_627: n_833  <= TRANSPORT NOT a_N1095_aNOT_aOUT  ;
delay_628: n_834  <= TRANSPORT a_N1094_aNOT_aOUT  ;
delay_629: n_835  <= TRANSPORT a_LC4_B2_aOUT  ;
and4_630: n_836 <=  n_837  AND n_838  AND n_839  AND n_840;
inv_631: n_837  <= TRANSPORT NOT a_N1096_aNOT_aOUT  ;
delay_632: n_838  <= TRANSPORT a_N1095_aNOT_aOUT  ;
inv_633: n_839  <= TRANSPORT NOT a_N1094_aNOT_aOUT  ;
delay_634: n_840  <= TRANSPORT a_LC4_B2_aOUT  ;
and4_635: n_841 <=  n_842  AND n_843  AND n_844  AND n_845;
delay_636: n_842  <= TRANSPORT a_N1096_aNOT_aOUT  ;
inv_637: n_843  <= TRANSPORT NOT a_N1095_aNOT_aOUT  ;
inv_638: n_844  <= TRANSPORT NOT a_N1094_aNOT_aOUT  ;
delay_639: n_845  <= TRANSPORT a_LC4_B2_aOUT  ;
and4_640: n_846 <=  n_847  AND n_848  AND n_849  AND n_850;
delay_641: n_847  <= TRANSPORT a_N1096_aNOT_aOUT  ;
delay_642: n_848  <= TRANSPORT a_N1095_aNOT_aOUT  ;
inv_643: n_849  <= TRANSPORT NOT a_N1094_aNOT_aOUT  ;
inv_644: n_850  <= TRANSPORT NOT a_LC4_B2_aOUT  ;
and4_645: n_851 <=  n_852  AND n_853  AND n_854  AND n_855;
inv_646: n_852  <= TRANSPORT NOT a_N1096_aNOT_aOUT  ;
inv_647: n_853  <= TRANSPORT NOT a_N1095_aNOT_aOUT  ;
inv_648: n_854  <= TRANSPORT NOT a_N1094_aNOT_aOUT  ;
inv_649: n_855  <= TRANSPORT NOT a_LC4_B2_aOUT  ;
and4_650: n_856 <=  n_857  AND n_858  AND n_859  AND n_860;
inv_651: n_857  <= TRANSPORT NOT a_N1096_aNOT_aOUT  ;
delay_652: n_858  <= TRANSPORT a_N1095_aNOT_aOUT  ;
delay_653: n_859  <= TRANSPORT a_N1094_aNOT_aOUT  ;
inv_654: n_860  <= TRANSPORT NOT a_LC4_B2_aOUT  ;
and4_655: n_861 <=  n_862  AND n_863  AND n_864  AND n_865;
delay_656: n_862  <= TRANSPORT a_N1096_aNOT_aOUT  ;
inv_657: n_863  <= TRANSPORT NOT a_N1095_aNOT_aOUT  ;
delay_658: n_864  <= TRANSPORT a_N1094_aNOT_aOUT  ;
inv_659: n_865  <= TRANSPORT NOT a_LC4_B2_aOUT  ;
and1_660: n_866 <=  gnd;
dff_661: DFF_a8251
    PORT MAP ( D => a_N868_aD, CLK => a_N868_aCLK, CLRN => a_N868_aCLRN, PRN => vcc,
          Q => a_N868_aQ);
delay_662: a_N868_aCLRN  <= TRANSPORT nRESET  ;
xor2_663: a_N868_aD <=  n_874  XOR n_886;
or3_664: n_874 <=  n_875  OR n_878  OR n_882;
and2_665: n_875 <=  n_876  AND n_877;
delay_666: n_876  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_667: n_877  <= TRANSPORT a_N868_aQ  ;
and3_668: n_878 <=  n_879  AND n_880  AND n_881;
inv_669: n_879  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_670: n_880  <= TRANSPORT a_LC8_B20_aOUT  ;
delay_671: n_881  <= TRANSPORT a_LC7_B2_aOUT  ;
and3_672: n_882 <=  n_883  AND n_884  AND n_885;
inv_673: n_883  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
inv_674: n_884  <= TRANSPORT NOT a_LC8_B20_aOUT  ;
inv_675: n_885  <= TRANSPORT NOT a_LC7_B2_aOUT  ;
and1_676: n_886 <=  gnd;
inv_677: n_887  <= TRANSPORT NOT nTXC  ;
filter_678: FILTER_a8251
    PORT MAP (IN1 => n_887, Y => a_N868_aCLK);
delay_679: a_LC5_B7_aOUT  <= TRANSPORT a_LC5_B7_aIN  ;
xor2_680: a_LC5_B7_aIN <=  n_891  XOR n_899;
or2_681: n_891 <=  n_892  OR n_896;
and2_682: n_892 <=  n_893  AND n_895;
inv_683: n_893  <= TRANSPORT NOT a_N1128_aNOT_aOUT  ;
delay_684: n_895  <= TRANSPORT a_STXRDY_aNOT_aQ  ;
and2_685: n_896 <=  n_897  AND n_898;
inv_686: n_897  <= TRANSPORT NOT a_N1128_aNOT_aOUT  ;
delay_687: n_898  <= TRANSPORT a_SMODE_OUT_F7_G_aQ  ;
and1_688: n_899 <=  gnd;
delay_689: a_N616_aOUT  <= TRANSPORT a_N616_aIN  ;
xor2_690: a_N616_aIN <=  n_902  XOR n_911;
or2_691: n_902 <=  n_903  OR n_907;
and2_692: n_903 <=  n_904  AND n_906;
inv_693: n_904  <= TRANSPORT NOT a_LC8_B4_aNOT_aOUT  ;
delay_694: n_906  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_695: n_907 <=  n_908  AND n_910;
inv_696: n_908  <= TRANSPORT NOT a_N80_aOUT  ;
delay_697: n_910  <= TRANSPORT a_LC5_B7_aOUT  ;
and1_698: n_911 <=  gnd;
delay_699: a_LC6_B7_aOUT  <= TRANSPORT a_LC6_B7_aIN  ;
xor2_700: a_LC6_B7_aIN <=  n_914  XOR n_922;
or2_701: n_914 <=  n_915  OR n_919;
and2_702: n_915 <=  n_916  AND n_918;
inv_703: n_916  <= TRANSPORT NOT a_N76_aNOT_aOUT  ;
delay_704: n_918  <= TRANSPORT a_N616_aOUT  ;
and1_705: n_919 <=  n_920;
inv_706: n_920  <= TRANSPORT NOT a_LC3_B7_aNOT_aOUT  ;
and1_707: n_922 <=  gnd;
delay_708: a_LC8_B7_aOUT  <= TRANSPORT a_LC8_B7_aIN  ;
xor2_709: a_LC8_B7_aIN <=  n_925  XOR n_935;
or3_710: n_925 <=  n_926  OR n_929  OR n_932;
and2_711: n_926 <=  n_927  AND n_928;
inv_712: n_927  <= TRANSPORT NOT a_N1128_aNOT_aOUT  ;
delay_713: n_928  <= TRANSPORT a_STXRDY_aNOT_aQ  ;
and2_714: n_929 <=  n_930  AND n_931;
delay_715: n_930  <= TRANSPORT a_N1107_aOUT  ;
inv_716: n_931  <= TRANSPORT NOT a_N1128_aNOT_aOUT  ;
and2_717: n_932 <=  n_933  AND n_934;
delay_718: n_933  <= TRANSPORT a_N80_aOUT  ;
delay_719: n_934  <= TRANSPORT a_N1128_aNOT_aOUT  ;
and1_720: n_935 <=  gnd;
dff_721: DFF_a8251
    PORT MAP ( D => a_N414_aD, CLK => a_N414_aCLK, CLRN => a_N414_aCLRN, PRN => vcc,
          Q => a_N414_aQ);
delay_722: a_N414_aCLRN  <= TRANSPORT nRESET  ;
xor2_723: a_N414_aD <=  n_942  XOR n_951;
or2_724: n_942 <=  n_943  OR n_947;
and3_725: n_943 <=  n_944  AND n_945  AND n_946;
delay_726: n_944  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_727: n_945  <= TRANSPORT a_LC6_B7_aOUT  ;
inv_728: n_946  <= TRANSPORT NOT a_N414_aQ  ;
and3_729: n_947 <=  n_948  AND n_949  AND n_950;
delay_730: n_948  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_731: n_949  <= TRANSPORT a_LC8_B7_aOUT  ;
delay_732: n_950  <= TRANSPORT a_N414_aQ  ;
and1_733: n_951 <=  gnd;
inv_734: n_952  <= TRANSPORT NOT nTXC  ;
filter_735: FILTER_a8251
    PORT MAP (IN1 => n_952, Y => a_N414_aCLK);
delay_736: a_LC2_B10_aOUT  <= TRANSPORT a_LC2_B10_aIN  ;
xor2_737: a_LC2_B10_aIN <=  n_956  XOR n_964;
or2_738: n_956 <=  n_957  OR n_961;
and2_739: n_957 <=  n_958  AND n_960;
inv_740: n_958  <= TRANSPORT NOT a_N1066_aNOT_aOUT  ;
delay_741: n_960  <= TRANSPORT a_N413_aQ  ;
and2_742: n_961 <=  n_962  AND n_963;
delay_743: n_962  <= TRANSPORT a_N80_aOUT  ;
delay_744: n_963  <= TRANSPORT a_N413_aQ  ;
and1_745: n_964 <=  gnd;
delay_746: a_LC2_B4_aOUT  <= TRANSPORT a_LC2_B4_aIN  ;
xor2_747: a_LC2_B4_aIN <=  n_967  XOR n_980;
or3_748: n_967 <=  n_968  OR n_973  OR n_977;
and2_749: n_968 <=  n_969  AND n_971;
inv_750: n_969  <= TRANSPORT NOT a_N1179_aNOT_aOUT  ;
inv_751: n_971  <= TRANSPORT NOT a_N394_aQ  ;
and2_752: n_973 <=  n_974  AND n_975;
inv_753: n_974  <= TRANSPORT NOT a_N1179_aNOT_aOUT  ;
delay_754: n_975  <= TRANSPORT a_LC1_B4_aNOT_aOUT  ;
and2_755: n_977 <=  n_978  AND n_979;
inv_756: n_978  <= TRANSPORT NOT a_N1179_aNOT_aOUT  ;
delay_757: n_979  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_758: n_980 <=  gnd;
dff_759: DFF_a8251
    PORT MAP ( D => a_N413_aD, CLK => a_N413_aCLK, CLRN => a_N413_aCLRN, PRN => vcc,
          Q => a_N413_aQ);
delay_760: a_N413_aCLRN  <= TRANSPORT nRESET  ;
xor2_761: a_N413_aD <=  n_987  XOR n_998;
or3_762: n_987 <=  n_988  OR n_991  OR n_994;
and2_763: n_988 <=  n_989  AND n_990;
delay_764: n_989  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_765: n_990  <= TRANSPORT a_LC2_B10_aOUT  ;
and2_766: n_991 <=  n_992  AND n_993;
delay_767: n_992  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_768: n_993  <= TRANSPORT a_LC2_B4_aOUT  ;
and2_769: n_994 <=  n_995  AND n_996;
delay_770: n_995  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_771: n_996  <= TRANSPORT NOT a_LC8_B10_aOUT  ;
and1_772: n_998 <=  gnd;
inv_773: n_999  <= TRANSPORT NOT nTXC  ;
filter_774: FILTER_a8251
    PORT MAP (IN1 => n_999, Y => a_N413_aCLK);
dff_775: DFF_a8251
    PORT MAP ( D => a_N1899_aD, CLK => a_N1899_aCLK, CLRN => a_N1899_aCLRN,
          PRN => vcc, Q => a_N1899_aQ);
delay_776: a_N1899_aCLRN  <= TRANSPORT nRESET  ;
xor2_777: a_N1899_aD <=  n_1008  XOR n_1012;
or1_778: n_1008 <=  n_1009;
and1_779: n_1009 <=  n_1010;
delay_780: n_1010  <= TRANSPORT a_N1900_aQ  ;
and1_781: n_1012 <=  gnd;
delay_782: n_1013  <= TRANSPORT nRXC  ;
filter_783: FILTER_a8251
    PORT MAP (IN1 => n_1013, Y => a_N1899_aCLK);
dff_784: DFF_a8251
    PORT MAP ( D => a_N1900_aD, CLK => a_N1900_aCLK, CLRN => a_N1900_aCLRN,
          PRN => vcc, Q => a_N1900_aQ);
delay_785: a_N1900_aCLRN  <= TRANSPORT nRESET  ;
xor2_786: a_N1900_aD <=  n_1021  XOR n_1027;
or1_787: n_1021 <=  n_1022;
and4_788: n_1022 <=  n_1023  AND n_1024  AND n_1025  AND n_1026;
delay_789: n_1023  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_790: n_1024  <= TRANSPORT a_N1754_aQ  ;
inv_791: n_1025  <= TRANSPORT NOT a_N1757_aQ  ;
inv_792: n_1026  <= TRANSPORT NOT a_N1756_aQ  ;
and1_793: n_1027 <=  gnd;
delay_794: n_1028  <= TRANSPORT nRXC  ;
filter_795: FILTER_a8251
    PORT MAP (IN1 => n_1028, Y => a_N1900_aCLK);
dff_796: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F0_G_aD, CLK => a_SCMND_OUT_F0_G_aCLK, CLRN => a_SCMND_OUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F0_G_aQ);
delay_797: a_SCMND_OUT_F0_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_798: a_SCMND_OUT_F0_G_aD <=  n_1037  XOR n_1046;
or2_799: n_1037 <=  n_1038  OR n_1042;
and3_800: n_1038 <=  n_1039  AND n_1040  AND n_1041;
delay_801: n_1039  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_802: n_1040  <= TRANSPORT NOT a_N701_aNOT_aOUT  ;
delay_803: n_1041  <= TRANSPORT a_SCMND_OUT_F0_G_aQ  ;
and3_804: n_1042 <=  n_1043  AND n_1044  AND n_1045;
delay_805: n_1043  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_806: n_1044  <= TRANSPORT a_N701_aNOT_aOUT  ;
delay_807: n_1045  <= TRANSPORT DIN(0)  ;
and1_808: n_1046 <=  gnd;
delay_809: n_1047  <= TRANSPORT CLK  ;
filter_810: FILTER_a8251
    PORT MAP (IN1 => n_1047, Y => a_SCMND_OUT_F0_G_aCLK);
dff_811: DFF_a8251
    PORT MAP ( D => a_SRXREG_F0_G_aD, CLK => a_SRXREG_F0_G_aCLK, CLRN => a_SRXREG_F0_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F0_G_aQ);
delay_812: a_SRXREG_F0_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_813: a_SRXREG_F0_G_aD <=  n_1056  XOR n_1068;
or2_814: n_1056 <=  n_1057  OR n_1063;
and3_815: n_1057 <=  n_1058  AND n_1060  AND n_1062;
inv_816: n_1058  <= TRANSPORT NOT a_N83_aOUT  ;
inv_817: n_1060  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_818: n_1062  <= TRANSPORT a_SRXREG_F0_G_aQ  ;
and3_819: n_1063 <=  n_1064  AND n_1065  AND n_1067;
inv_820: n_1064  <= TRANSPORT NOT a_N83_aOUT  ;
delay_821: n_1065  <= TRANSPORT a_N1100_aNOT_aOUT  ;
delay_822: n_1067  <= TRANSPORT a_N79_aNOT_aOUT  ;
and1_823: n_1068 <=  gnd;
delay_824: n_1069  <= TRANSPORT nRXC  ;
filter_825: FILTER_a8251
    PORT MAP (IN1 => n_1069, Y => a_SRXREG_F0_G_aCLK);
dff_826: DFF_a8251
    PORT MAP ( D => a_SRXREG_F1_G_aD, CLK => a_SRXREG_F1_G_aCLK, CLRN => a_SRXREG_F1_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F1_G_aQ);
delay_827: a_SRXREG_F1_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_828: a_SRXREG_F1_G_aD <=  n_1078  XOR n_1088;
or2_829: n_1078 <=  n_1079  OR n_1083;
and3_830: n_1079 <=  n_1080  AND n_1081  AND n_1082;
inv_831: n_1080  <= TRANSPORT NOT a_N83_aOUT  ;
inv_832: n_1081  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_833: n_1082  <= TRANSPORT a_SRXREG_F1_G_aQ  ;
and3_834: n_1083 <=  n_1084  AND n_1085  AND n_1087;
inv_835: n_1084  <= TRANSPORT NOT a_N83_aOUT  ;
delay_836: n_1085  <= TRANSPORT a_N1101_aNOT_aOUT  ;
delay_837: n_1087  <= TRANSPORT a_N79_aNOT_aOUT  ;
and1_838: n_1088 <=  gnd;
delay_839: n_1089  <= TRANSPORT nRXC  ;
filter_840: FILTER_a8251
    PORT MAP (IN1 => n_1089, Y => a_SRXREG_F1_G_aCLK);
dff_841: DFF_a8251
    PORT MAP ( D => a_SRXREG_F2_G_aD, CLK => a_SRXREG_F2_G_aCLK, CLRN => a_SRXREG_F2_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F2_G_aQ);
delay_842: a_SRXREG_F2_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_843: a_SRXREG_F2_G_aD <=  n_1098  XOR n_1109;
or2_844: n_1098 <=  n_1099  OR n_1104;
and3_845: n_1099 <=  n_1100  AND n_1101  AND n_1103;
inv_846: n_1100  <= TRANSPORT NOT a_N83_aOUT  ;
inv_847: n_1101  <= TRANSPORT NOT a_N134_aNOT_aOUT  ;
delay_848: n_1103  <= TRANSPORT a_SRXREG_F2_G_aQ  ;
and3_849: n_1104 <=  n_1105  AND n_1106  AND n_1108;
inv_850: n_1105  <= TRANSPORT NOT a_N83_aOUT  ;
delay_851: n_1106  <= TRANSPORT a_N1102_aNOT_aOUT  ;
delay_852: n_1108  <= TRANSPORT a_N134_aNOT_aOUT  ;
and1_853: n_1109 <=  gnd;
delay_854: n_1110  <= TRANSPORT nRXC  ;
filter_855: FILTER_a8251
    PORT MAP (IN1 => n_1110, Y => a_SRXREG_F2_G_aCLK);
dff_856: DFF_a8251
    PORT MAP ( D => a_SRXREG_F3_G_aD, CLK => a_SRXREG_F3_G_aCLK, CLRN => a_SRXREG_F3_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F3_G_aQ);
delay_857: a_SRXREG_F3_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_858: a_SRXREG_F3_G_aD <=  n_1119  XOR n_1129;
or2_859: n_1119 <=  n_1120  OR n_1125;
and3_860: n_1120 <=  n_1121  AND n_1122  AND n_1124;
inv_861: n_1121  <= TRANSPORT NOT a_N83_aOUT  ;
delay_862: n_1122  <= TRANSPORT a_N1103_aNOT_aOUT  ;
delay_863: n_1124  <= TRANSPORT a_N79_aNOT_aOUT  ;
and3_864: n_1125 <=  n_1126  AND n_1127  AND n_1128;
inv_865: n_1126  <= TRANSPORT NOT a_N83_aOUT  ;
inv_866: n_1127  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_867: n_1128  <= TRANSPORT a_SRXREG_F3_G_aQ  ;
and1_868: n_1129 <=  gnd;
delay_869: n_1130  <= TRANSPORT nRXC  ;
filter_870: FILTER_a8251
    PORT MAP (IN1 => n_1130, Y => a_SRXREG_F3_G_aCLK);
delay_871: a_LC7_A11_aOUT  <= TRANSPORT a_LC7_A11_aIN  ;
xor2_872: a_LC7_A11_aIN <=  n_1134  XOR n_1176;
or8_873: n_1134 <=  n_1135  OR n_1141  OR n_1146  OR n_1151  OR n_1156  OR n_1161
           OR n_1166  OR n_1171;
and4_874: n_1135 <=  n_1136  AND n_1137  AND n_1138  AND n_1139;
delay_875: n_1136  <= TRANSPORT a_N1102_aNOT_aOUT  ;
inv_876: n_1137  <= TRANSPORT NOT a_N1101_aNOT_aOUT  ;
delay_877: n_1138  <= TRANSPORT a_N1100_aNOT_aOUT  ;
delay_878: n_1139  <= TRANSPORT a_N1106_aNOT_aOUT  ;
and4_879: n_1141 <=  n_1142  AND n_1143  AND n_1144  AND n_1145;
delay_880: n_1142  <= TRANSPORT a_N1102_aNOT_aOUT  ;
delay_881: n_1143  <= TRANSPORT a_N1101_aNOT_aOUT  ;
delay_882: n_1144  <= TRANSPORT a_N1100_aNOT_aOUT  ;
inv_883: n_1145  <= TRANSPORT NOT a_N1106_aNOT_aOUT  ;
and4_884: n_1146 <=  n_1147  AND n_1148  AND n_1149  AND n_1150;
delay_885: n_1147  <= TRANSPORT a_N1102_aNOT_aOUT  ;
inv_886: n_1148  <= TRANSPORT NOT a_N1101_aNOT_aOUT  ;
inv_887: n_1149  <= TRANSPORT NOT a_N1100_aNOT_aOUT  ;
inv_888: n_1150  <= TRANSPORT NOT a_N1106_aNOT_aOUT  ;
and4_889: n_1151 <=  n_1152  AND n_1153  AND n_1154  AND n_1155;
delay_890: n_1152  <= TRANSPORT a_N1102_aNOT_aOUT  ;
delay_891: n_1153  <= TRANSPORT a_N1101_aNOT_aOUT  ;
inv_892: n_1154  <= TRANSPORT NOT a_N1100_aNOT_aOUT  ;
delay_893: n_1155  <= TRANSPORT a_N1106_aNOT_aOUT  ;
and4_894: n_1156 <=  n_1157  AND n_1158  AND n_1159  AND n_1160;
inv_895: n_1157  <= TRANSPORT NOT a_N1102_aNOT_aOUT  ;
inv_896: n_1158  <= TRANSPORT NOT a_N1101_aNOT_aOUT  ;
inv_897: n_1159  <= TRANSPORT NOT a_N1100_aNOT_aOUT  ;
delay_898: n_1160  <= TRANSPORT a_N1106_aNOT_aOUT  ;
and4_899: n_1161 <=  n_1162  AND n_1163  AND n_1164  AND n_1165;
inv_900: n_1162  <= TRANSPORT NOT a_N1102_aNOT_aOUT  ;
delay_901: n_1163  <= TRANSPORT a_N1101_aNOT_aOUT  ;
inv_902: n_1164  <= TRANSPORT NOT a_N1100_aNOT_aOUT  ;
inv_903: n_1165  <= TRANSPORT NOT a_N1106_aNOT_aOUT  ;
and4_904: n_1166 <=  n_1167  AND n_1168  AND n_1169  AND n_1170;
inv_905: n_1167  <= TRANSPORT NOT a_N1102_aNOT_aOUT  ;
inv_906: n_1168  <= TRANSPORT NOT a_N1101_aNOT_aOUT  ;
delay_907: n_1169  <= TRANSPORT a_N1100_aNOT_aOUT  ;
inv_908: n_1170  <= TRANSPORT NOT a_N1106_aNOT_aOUT  ;
and4_909: n_1171 <=  n_1172  AND n_1173  AND n_1174  AND n_1175;
inv_910: n_1172  <= TRANSPORT NOT a_N1102_aNOT_aOUT  ;
delay_911: n_1173  <= TRANSPORT a_N1101_aNOT_aOUT  ;
delay_912: n_1174  <= TRANSPORT a_N1100_aNOT_aOUT  ;
delay_913: n_1175  <= TRANSPORT a_N1106_aNOT_aOUT  ;
and1_914: n_1176 <=  gnd;
delay_915: a_LC1_A11_aOUT  <= TRANSPORT a_LC1_A11_aIN  ;
xor2_916: a_LC1_A11_aIN <=  n_1179  XOR n_1222;
or8_917: n_1179 <=  n_1180  OR n_1187  OR n_1192  OR n_1197  OR n_1202  OR n_1207
           OR n_1212  OR n_1217;
and4_918: n_1180 <=  n_1181  AND n_1183  AND n_1184  AND n_1186;
delay_919: n_1181  <= TRANSPORT a_N1105_aNOT_aOUT  ;
delay_920: n_1183  <= TRANSPORT a_N1103_aNOT_aOUT  ;
delay_921: n_1184  <= TRANSPORT a_N96_aOUT  ;
delay_922: n_1186  <= TRANSPORT a_LC7_A11_aOUT  ;
and4_923: n_1187 <=  n_1188  AND n_1189  AND n_1190  AND n_1191;
inv_924: n_1188  <= TRANSPORT NOT a_N1105_aNOT_aOUT  ;
delay_925: n_1189  <= TRANSPORT a_N1103_aNOT_aOUT  ;
inv_926: n_1190  <= TRANSPORT NOT a_N96_aOUT  ;
delay_927: n_1191  <= TRANSPORT a_LC7_A11_aOUT  ;
and4_928: n_1192 <=  n_1193  AND n_1194  AND n_1195  AND n_1196;
delay_929: n_1193  <= TRANSPORT a_N1105_aNOT_aOUT  ;
inv_930: n_1194  <= TRANSPORT NOT a_N1103_aNOT_aOUT  ;
inv_931: n_1195  <= TRANSPORT NOT a_N96_aOUT  ;
delay_932: n_1196  <= TRANSPORT a_LC7_A11_aOUT  ;
and4_933: n_1197 <=  n_1198  AND n_1199  AND n_1200  AND n_1201;
inv_934: n_1198  <= TRANSPORT NOT a_N1105_aNOT_aOUT  ;
inv_935: n_1199  <= TRANSPORT NOT a_N1103_aNOT_aOUT  ;
delay_936: n_1200  <= TRANSPORT a_N96_aOUT  ;
delay_937: n_1201  <= TRANSPORT a_LC7_A11_aOUT  ;
and4_938: n_1202 <=  n_1203  AND n_1204  AND n_1205  AND n_1206;
delay_939: n_1203  <= TRANSPORT a_N1105_aNOT_aOUT  ;
inv_940: n_1204  <= TRANSPORT NOT a_N1103_aNOT_aOUT  ;
delay_941: n_1205  <= TRANSPORT a_N96_aOUT  ;
inv_942: n_1206  <= TRANSPORT NOT a_LC7_A11_aOUT  ;
and4_943: n_1207 <=  n_1208  AND n_1209  AND n_1210  AND n_1211;
inv_944: n_1208  <= TRANSPORT NOT a_N1105_aNOT_aOUT  ;
inv_945: n_1209  <= TRANSPORT NOT a_N1103_aNOT_aOUT  ;
inv_946: n_1210  <= TRANSPORT NOT a_N96_aOUT  ;
inv_947: n_1211  <= TRANSPORT NOT a_LC7_A11_aOUT  ;
and4_948: n_1212 <=  n_1213  AND n_1214  AND n_1215  AND n_1216;
delay_949: n_1213  <= TRANSPORT a_N1105_aNOT_aOUT  ;
delay_950: n_1214  <= TRANSPORT a_N1103_aNOT_aOUT  ;
inv_951: n_1215  <= TRANSPORT NOT a_N96_aOUT  ;
inv_952: n_1216  <= TRANSPORT NOT a_LC7_A11_aOUT  ;
and4_953: n_1217 <=  n_1218  AND n_1219  AND n_1220  AND n_1221;
inv_954: n_1218  <= TRANSPORT NOT a_N1105_aNOT_aOUT  ;
delay_955: n_1219  <= TRANSPORT a_N1103_aNOT_aOUT  ;
delay_956: n_1220  <= TRANSPORT a_N96_aOUT  ;
inv_957: n_1221  <= TRANSPORT NOT a_LC7_A11_aOUT  ;
and1_958: n_1222 <=  gnd;
delay_959: a_N552_aNOT_aOUT  <= TRANSPORT a_N552_aNOT_aIN  ;
xor2_960: a_N552_aNOT_aIN <=  n_1225  XOR n_1240;
or4_961: n_1225 <=  n_1226  OR n_1230  OR n_1233  OR n_1237;
and2_962: n_1226 <=  n_1227  AND n_1229;
delay_963: n_1227  <= TRANSPORT a_N1104_aNOT_aOUT  ;
delay_964: n_1229  <= TRANSPORT a_LC1_A11_aOUT  ;
and2_965: n_1230 <=  n_1231  AND n_1232;
inv_966: n_1231  <= TRANSPORT NOT a_N1104_aNOT_aOUT  ;
inv_967: n_1232  <= TRANSPORT NOT a_LC1_A11_aOUT  ;
and2_968: n_1233 <=  n_1234  AND n_1236;
inv_969: n_1234  <= TRANSPORT NOT a_N1998_aQ  ;
inv_970: n_1236  <= TRANSPORT NOT a_SMODE_OUT_F5_G_aQ  ;
and2_971: n_1237 <=  n_1238  AND n_1239;
delay_972: n_1238  <= TRANSPORT a_N1998_aQ  ;
delay_973: n_1239  <= TRANSPORT a_SMODE_OUT_F5_G_aQ  ;
and1_974: n_1240 <=  gnd;
delay_975: a_N551_aNOT_aOUT  <= TRANSPORT a_N551_aNOT_aIN  ;
xor2_976: a_N551_aNOT_aIN <=  n_1243  XOR n_1256;
or4_977: n_1243 <=  n_1244  OR n_1247  OR n_1250  OR n_1253;
and2_978: n_1244 <=  n_1245  AND n_1246;
inv_979: n_1245  <= TRANSPORT NOT a_N1104_aNOT_aOUT  ;
delay_980: n_1246  <= TRANSPORT a_LC1_A11_aOUT  ;
and2_981: n_1247 <=  n_1248  AND n_1249;
delay_982: n_1248  <= TRANSPORT a_N1104_aNOT_aOUT  ;
inv_983: n_1249  <= TRANSPORT NOT a_LC1_A11_aOUT  ;
and2_984: n_1250 <=  n_1251  AND n_1252;
inv_985: n_1251  <= TRANSPORT NOT a_N1998_aQ  ;
delay_986: n_1252  <= TRANSPORT a_SMODE_OUT_F5_G_aQ  ;
and2_987: n_1253 <=  n_1254  AND n_1255;
delay_988: n_1254  <= TRANSPORT a_N1998_aQ  ;
inv_989: n_1255  <= TRANSPORT NOT a_SMODE_OUT_F5_G_aQ  ;
and1_990: n_1256 <=  gnd;
delay_991: a_LC2_C6_aOUT  <= TRANSPORT a_LC2_C6_aIN  ;
xor2_992: a_LC2_C6_aIN <=  n_1259  XOR n_1265;
or1_993: n_1259 <=  n_1260;
and4_994: n_1260 <=  n_1261  AND n_1262  AND n_1263  AND n_1264;
inv_995: n_1261  <= TRANSPORT NOT a_N83_aOUT  ;
delay_996: n_1262  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
delay_997: n_1263  <= TRANSPORT a_N552_aNOT_aOUT  ;
delay_998: n_1264  <= TRANSPORT a_N551_aNOT_aOUT  ;
and1_999: n_1265 <=  gnd;
delay_1000: a_LC5_C21_aOUT  <= TRANSPORT a_LC5_C21_aIN  ;
xor2_1001: a_LC5_C21_aIN <=  n_1268  XOR n_1277;
or2_1002: n_1268 <=  n_1269  OR n_1274;
and3_1003: n_1269 <=  n_1270  AND n_1271  AND n_1272;
inv_1004: n_1270  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1005: n_1271  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_1006: n_1272  <= TRANSPORT pe_aQ  ;
and2_1007: n_1274 <=  n_1275  AND n_1276;
delay_1008: n_1275  <= TRANSPORT a_N79_aNOT_aOUT  ;
delay_1009: n_1276  <= TRANSPORT a_LC2_C6_aOUT  ;
and1_1010: n_1277 <=  gnd;
dff_1011: DFF_a8251
    PORT MAP ( D => pe_aD, CLK => pe_aCLK, CLRN => pe_aCLRN, PRN => vcc, Q => pe_aQ);
delay_1012: pe_aCLRN  <= TRANSPORT nRESET  ;
xor2_1013: pe_aD <=  n_1284  XOR n_1291;
or2_1014: n_1284 <=  n_1285  OR n_1288;
and2_1015: n_1285 <=  n_1286  AND n_1287;
inv_1016: n_1286  <= TRANSPORT NOT a_N1898_aQ  ;
delay_1017: n_1287  <= TRANSPORT a_LC5_C21_aOUT  ;
and2_1018: n_1288 <=  n_1289  AND n_1290;
delay_1019: n_1289  <= TRANSPORT a_N1897_aQ  ;
delay_1020: n_1290  <= TRANSPORT a_LC5_C21_aOUT  ;
and1_1021: n_1291 <=  gnd;
delay_1022: n_1292  <= TRANSPORT nRXC  ;
filter_1023: FILTER_a8251
    PORT MAP (IN1 => n_1292, Y => pe_aCLK);
dff_1024: DFF_a8251
    PORT MAP ( D => a_SRXREG_F4_G_aD, CLK => a_SRXREG_F4_G_aCLK, CLRN => a_SRXREG_F4_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F4_G_aQ);
delay_1025: a_SRXREG_F4_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1026: a_SRXREG_F4_G_aD <=  n_1301  XOR n_1310;
or2_1027: n_1301 <=  n_1302  OR n_1306;
and3_1028: n_1302 <=  n_1303  AND n_1304  AND n_1305;
inv_1029: n_1303  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1030: n_1304  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_1031: n_1305  <= TRANSPORT a_SRXREG_F4_G_aQ  ;
and3_1032: n_1306 <=  n_1307  AND n_1308  AND n_1309;
inv_1033: n_1307  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1034: n_1308  <= TRANSPORT a_N1104_aNOT_aOUT  ;
delay_1035: n_1309  <= TRANSPORT a_N79_aNOT_aOUT  ;
and1_1036: n_1310 <=  gnd;
delay_1037: n_1311  <= TRANSPORT nRXC  ;
filter_1038: FILTER_a8251
    PORT MAP (IN1 => n_1311, Y => a_SRXREG_F4_G_aCLK);
delay_1039: a_N325_aNOT_aOUT  <= TRANSPORT a_N325_aNOT_aIN  ;
xor2_1040: a_N325_aNOT_aIN <=  n_1315  XOR n_1329;
or2_1041: n_1315 <=  n_1316  OR n_1325;
and4_1042: n_1316 <=  n_1317  AND n_1319  AND n_1321  AND n_1323;
inv_1043: n_1317  <= TRANSPORT NOT a_N1163_aNOT_aOUT  ;
delay_1044: n_1319  <= TRANSPORT a_N59_aQ  ;
inv_1045: n_1321  <= TRANSPORT NOT a_N62_aQ  ;
inv_1046: n_1323  <= TRANSPORT NOT a_N61_aQ  ;
and3_1047: n_1325 <=  n_1326  AND n_1327  AND n_1328;
inv_1048: n_1326  <= TRANSPORT NOT a_N1163_aNOT_aOUT  ;
delay_1049: n_1327  <= TRANSPORT a_N62_aQ  ;
delay_1050: n_1328  <= TRANSPORT a_N61_aQ  ;
and1_1051: n_1329 <=  gnd;
delay_1052: a_N329_aNOT_aOUT  <= TRANSPORT a_N329_aNOT_aIN  ;
xor2_1053: a_N329_aNOT_aIN <=  n_1332  XOR n_1342;
or1_1054: n_1332 <=  n_1333;
and4_1055: n_1333 <=  n_1334  AND n_1336  AND n_1338  AND n_1340;
delay_1056: n_1334  <= TRANSPORT a_N1183_aNOT_aOUT  ;
delay_1057: n_1336  <= TRANSPORT a_N1145_aOUT  ;
delay_1058: n_1338  <= TRANSPORT a_N64_aQ  ;
inv_1059: n_1340  <= TRANSPORT NOT a_N63_aQ  ;
and1_1060: n_1342 <=  gnd;
delay_1061: a_LC3_D3_aOUT  <= TRANSPORT a_LC3_D3_aIN  ;
xor2_1062: a_LC3_D3_aIN <=  n_1345  XOR n_1356;
or3_1063: n_1345 <=  n_1346  OR n_1349  OR n_1352;
and2_1064: n_1346 <=  n_1347  AND n_1348;
delay_1065: n_1347  <= TRANSPORT a_N325_aNOT_aOUT  ;
delay_1066: n_1348  <= TRANSPORT a_SRXRDY_aQ  ;
and2_1067: n_1349 <=  n_1350  AND n_1351;
delay_1068: n_1350  <= TRANSPORT a_N329_aNOT_aOUT  ;
delay_1069: n_1351  <= TRANSPORT a_SRXRDY_aQ  ;
and2_1070: n_1352 <=  n_1353  AND n_1355;
delay_1071: n_1353  <= TRANSPORT a_LC6_D4_aOUT  ;
delay_1072: n_1355  <= TRANSPORT a_SRXRDY_aQ  ;
and1_1073: n_1356 <=  gnd;
dff_1074: DFF_a8251
    PORT MAP ( D => oe_aD, CLK => oe_aCLK, CLRN => oe_aCLRN, PRN => vcc, Q => oe_aQ);
delay_1075: oe_aCLRN  <= TRANSPORT nRESET  ;
xor2_1076: oe_aD <=  n_1364  XOR n_1373;
or2_1077: n_1364 <=  n_1365  OR n_1369;
and3_1078: n_1365 <=  n_1366  AND n_1367  AND n_1368;
inv_1079: n_1366  <= TRANSPORT NOT a_N134_aNOT_aOUT  ;
inv_1080: n_1367  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_1081: n_1368  <= TRANSPORT oe_aQ  ;
and3_1082: n_1369 <=  n_1370  AND n_1371  AND n_1372;
delay_1083: n_1370  <= TRANSPORT a_N134_aNOT_aOUT  ;
inv_1084: n_1371  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_1085: n_1372  <= TRANSPORT a_LC3_D3_aOUT  ;
and1_1086: n_1373 <=  gnd;
delay_1087: n_1374  <= TRANSPORT nRXC  ;
filter_1088: FILTER_a8251
    PORT MAP (IN1 => n_1374, Y => oe_aCLK);
delay_1089: a_LC4_D20_aOUT  <= TRANSPORT a_LC4_D20_aIN  ;
xor2_1090: a_LC4_D20_aIN <=  n_1378  XOR n_1387;
or2_1091: n_1378 <=  n_1379  OR n_1383;
and3_1092: n_1379 <=  n_1380  AND n_1381  AND n_1382;
inv_1093: n_1380  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1094: n_1381  <= TRANSPORT a_N1105_aNOT_aOUT  ;
delay_1095: n_1382  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and3_1096: n_1383 <=  n_1384  AND n_1385  AND n_1386;
inv_1097: n_1384  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1098: n_1385  <= TRANSPORT a_N1105_aNOT_aOUT  ;
delay_1099: n_1386  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_1100: n_1387 <=  gnd;
dff_1101: DFF_a8251
    PORT MAP ( D => a_SRXREG_F5_G_aD, CLK => a_SRXREG_F5_G_aCLK, CLRN => a_SRXREG_F5_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F5_G_aQ);
delay_1102: a_SRXREG_F5_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1103: a_SRXREG_F5_G_aD <=  n_1395  XOR n_1404;
or2_1104: n_1395 <=  n_1396  OR n_1400;
and3_1105: n_1396 <=  n_1397  AND n_1398  AND n_1399;
inv_1106: n_1397  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1107: n_1398  <= TRANSPORT a_N79_aNOT_aOUT  ;
delay_1108: n_1399  <= TRANSPORT a_LC4_D20_aOUT  ;
and3_1109: n_1400 <=  n_1401  AND n_1402  AND n_1403;
inv_1110: n_1401  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1111: n_1402  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_1112: n_1403  <= TRANSPORT a_SRXREG_F5_G_aQ  ;
and1_1113: n_1404 <=  gnd;
delay_1114: n_1405  <= TRANSPORT nRXC  ;
filter_1115: FILTER_a8251
    PORT MAP (IN1 => n_1405, Y => a_SRXREG_F5_G_aCLK);
delay_1116: a_N708_aNOT_aOUT  <= TRANSPORT a_N708_aNOT_aIN  ;
xor2_1117: a_N708_aNOT_aIN <=  n_1409  XOR n_1414;
or1_1118: n_1409 <=  n_1410;
and3_1119: n_1410 <=  n_1411  AND n_1412  AND n_1413;
delay_1120: n_1411  <= TRANSPORT a_N1145_aOUT  ;
delay_1121: n_1412  <= TRANSPORT a_N64_aQ  ;
inv_1122: n_1413  <= TRANSPORT NOT a_N63_aQ  ;
and1_1123: n_1414 <=  gnd;
delay_1124: a_N707_aNOT_aOUT  <= TRANSPORT a_N707_aNOT_aIN  ;
xor2_1125: a_N707_aNOT_aIN <=  n_1417  XOR n_1428;
or2_1126: n_1417 <=  n_1418  OR n_1423;
and3_1127: n_1418 <=  n_1419  AND n_1420  AND n_1422;
inv_1128: n_1419  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1129: n_1420  <= TRANSPORT NOT RXD  ;
delay_1130: n_1422  <= TRANSPORT a_N708_aNOT_aOUT  ;
and3_1131: n_1423 <=  n_1424  AND n_1425  AND n_1427;
inv_1132: n_1424  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1133: n_1425  <= TRANSPORT a_N141_aNOT_aOUT  ;
inv_1134: n_1427  <= TRANSPORT NOT RXD  ;
and1_1135: n_1428 <=  gnd;
dff_1136: DFF_a8251
    PORT MAP ( D => fe_aD, CLK => fe_aCLK, CLRN => fe_aCLRN, PRN => vcc, Q => fe_aQ);
delay_1137: fe_aCLRN  <= TRANSPORT nRESET  ;
xor2_1138: fe_aD <=  n_1436  XOR n_1443;
or2_1139: n_1436 <=  n_1437  OR n_1440;
and2_1140: n_1437 <=  n_1438  AND n_1439;
inv_1141: n_1438  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_1142: n_1439  <= TRANSPORT fe_aQ  ;
and2_1143: n_1440 <=  n_1441  AND n_1442;
inv_1144: n_1441  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_1145: n_1442  <= TRANSPORT a_N707_aNOT_aOUT  ;
and1_1146: n_1443 <=  gnd;
delay_1147: n_1444  <= TRANSPORT nRXC  ;
filter_1148: FILTER_a8251
    PORT MAP (IN1 => n_1444, Y => fe_aCLK);
delay_1149: a_LC1_C6_aOUT  <= TRANSPORT a_LC1_C6_aIN  ;
xor2_1150: a_LC1_C6_aIN <=  n_1448  XOR n_1452;
or1_1151: n_1448 <=  n_1449;
and2_1152: n_1449 <=  n_1450  AND n_1451;
delay_1153: n_1450  <= TRANSPORT a_N1106_aNOT_aOUT  ;
delay_1154: n_1451  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_1155: n_1452 <=  gnd;
dff_1156: DFF_a8251
    PORT MAP ( D => a_SRXREG_F6_G_aD, CLK => a_SRXREG_F6_G_aCLK, CLRN => a_SRXREG_F6_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F6_G_aQ);
delay_1157: a_SRXREG_F6_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1158: a_SRXREG_F6_G_aD <=  n_1460  XOR n_1469;
or2_1159: n_1460 <=  n_1461  OR n_1465;
and3_1160: n_1461 <=  n_1462  AND n_1463  AND n_1464;
inv_1161: n_1462  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1162: n_1463  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_1163: n_1464  <= TRANSPORT a_SRXREG_F6_G_aQ  ;
and3_1164: n_1465 <=  n_1466  AND n_1467  AND n_1468;
inv_1165: n_1466  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1166: n_1467  <= TRANSPORT a_N79_aNOT_aOUT  ;
delay_1167: n_1468  <= TRANSPORT a_LC1_C6_aOUT  ;
and1_1168: n_1469 <=  gnd;
delay_1169: n_1470  <= TRANSPORT nRXC  ;
filter_1170: FILTER_a8251
    PORT MAP (IN1 => n_1470, Y => a_SRXREG_F6_G_aCLK);
dff_1171: DFF_a8251
    PORT MAP ( D => a_SRXREG_F7_G_aD, CLK => a_SRXREG_F7_G_aCLK, CLRN => a_SRXREG_F7_G_aCLRN,
          PRN => vcc, Q => a_SRXREG_F7_G_aQ);
delay_1172: a_SRXREG_F7_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1173: a_SRXREG_F7_G_aD <=  n_1479  XOR n_1488;
or2_1174: n_1479 <=  n_1480  OR n_1484;
and3_1175: n_1480 <=  n_1481  AND n_1482  AND n_1483;
inv_1176: n_1481  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1177: n_1482  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_1178: n_1483  <= TRANSPORT a_SRXREG_F7_G_aQ  ;
and3_1179: n_1484 <=  n_1485  AND n_1486  AND n_1487;
inv_1180: n_1485  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1181: n_1486  <= TRANSPORT a_N96_aOUT  ;
delay_1182: n_1487  <= TRANSPORT a_N79_aNOT_aOUT  ;
and1_1183: n_1488 <=  gnd;
delay_1184: n_1489  <= TRANSPORT nRXC  ;
filter_1185: FILTER_a8251
    PORT MAP (IN1 => n_1489, Y => a_SRXREG_F7_G_aCLK);
delay_1186: a_LC4_C7_aOUT  <= TRANSPORT a_LC4_C7_aIN  ;
xor2_1187: a_LC4_C7_aIN <=  n_1493  XOR n_1504;
or2_1188: n_1493 <=  n_1494  OR n_1500;
and3_1189: n_1494 <=  n_1495  AND n_1497  AND n_1498;
inv_1190: n_1495  <= TRANSPORT NOT a_N1120_aNOT_aOUT  ;
inv_1191: n_1497  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_1192: n_1498  <= TRANSPORT a_SCMND_OUT_F3_G_aQ  ;
and2_1193: n_1500 <=  n_1501  AND n_1503;
delay_1194: n_1501  <= TRANSPORT a_N613_aOUT  ;
delay_1195: n_1503  <= TRANSPORT a_SCMND_OUT_F3_G_aQ  ;
and1_1196: n_1504 <=  gnd;
dff_1197: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F3_G_aD, CLK => a_SCMND_OUT_F3_G_aCLK, CLRN => a_SCMND_OUT_F3_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F3_G_aQ);
delay_1198: a_SCMND_OUT_F3_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1199: a_SCMND_OUT_F3_G_aD <=  n_1511  XOR n_1519;
or2_1200: n_1511 <=  n_1512  OR n_1515;
and2_1201: n_1512 <=  n_1513  AND n_1514;
delay_1202: n_1513  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1203: n_1514  <= TRANSPORT a_LC4_C7_aOUT  ;
and3_1204: n_1515 <=  n_1516  AND n_1517  AND n_1518;
delay_1205: n_1516  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1206: n_1517  <= TRANSPORT a_N701_aNOT_aOUT  ;
delay_1207: n_1518  <= TRANSPORT DIN(3)  ;
and1_1208: n_1519 <=  gnd;
delay_1209: n_1520  <= TRANSPORT CLK  ;
filter_1210: FILTER_a8251
    PORT MAP (IN1 => n_1520, Y => a_SCMND_OUT_F3_G_aCLK);
delay_1211: a_LC2_C4_aOUT  <= TRANSPORT a_LC2_C4_aIN  ;
xor2_1212: a_LC2_C4_aIN <=  n_1524  XOR n_1530;
or1_1213: n_1524 <=  n_1525;
and4_1214: n_1525 <=  n_1526  AND n_1527  AND n_1528  AND n_1529;
delay_1215: n_1526  <= TRANSPORT a_LC1_C2_aOUT  ;
delay_1216: n_1527  <= TRANSPORT a_N1804_aQ  ;
inv_1217: n_1528  <= TRANSPORT NOT a_N1807_aQ  ;
delay_1218: n_1529  <= TRANSPORT DIN(0)  ;
and1_1219: n_1530 <=  gnd;
dff_1220: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F0_G_aD, CLK => a_SMODE_OUT_F0_G_aCLK, CLRN => a_SMODE_OUT_F0_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F0_G_aQ);
delay_1221: a_SMODE_OUT_F0_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1222: a_SMODE_OUT_F0_G_aD <=  n_1537  XOR n_1545;
or2_1223: n_1537 <=  n_1538  OR n_1541;
and2_1224: n_1538 <=  n_1539  AND n_1540;
delay_1225: n_1539  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1226: n_1540  <= TRANSPORT a_LC2_C4_aOUT  ;
and3_1227: n_1541 <=  n_1542  AND n_1543  AND n_1544;
delay_1228: n_1542  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1229: n_1543  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_1230: n_1544  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and1_1231: n_1545 <=  gnd;
delay_1232: n_1546  <= TRANSPORT CLK  ;
filter_1233: FILTER_a8251
    PORT MAP (IN1 => n_1546, Y => a_SMODE_OUT_F0_G_aCLK);
delay_1234: a_LC6_C4_aOUT  <= TRANSPORT a_LC6_C4_aIN  ;
xor2_1235: a_LC6_C4_aIN <=  n_1550  XOR n_1557;
or1_1236: n_1550 <=  n_1551;
and4_1237: n_1551 <=  n_1552  AND n_1553  AND n_1554  AND n_1555;
inv_1238: n_1552  <= TRANSPORT NOT a_N1123_aNOT_aOUT  ;
delay_1239: n_1553  <= TRANSPORT a_N1804_aQ  ;
inv_1240: n_1554  <= TRANSPORT NOT a_N1807_aQ  ;
delay_1241: n_1555  <= TRANSPORT DIN(1)  ;
and1_1242: n_1557 <=  gnd;
dff_1243: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F1_G_aD, CLK => a_SMODE_OUT_F1_G_aCLK, CLRN => a_SMODE_OUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F1_G_aQ);
delay_1244: a_SMODE_OUT_F1_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1245: a_SMODE_OUT_F1_G_aD <=  n_1564  XOR n_1572;
or2_1246: n_1564 <=  n_1565  OR n_1569;
and3_1247: n_1565 <=  n_1566  AND n_1567  AND n_1568;
delay_1248: n_1566  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1249: n_1567  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_1250: n_1568  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and2_1251: n_1569 <=  n_1570  AND n_1571;
delay_1252: n_1570  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1253: n_1571  <= TRANSPORT a_LC6_C4_aOUT  ;
and1_1254: n_1572 <=  gnd;
delay_1255: n_1573  <= TRANSPORT CLK  ;
filter_1256: FILTER_a8251
    PORT MAP (IN1 => n_1573, Y => a_SMODE_OUT_F1_G_aCLK);
delay_1257: a_SNEN_aNOT_aOUT  <= TRANSPORT a_SNEN_aNOT_aIN  ;
xor2_1258: a_SNEN_aNOT_aIN <=  n_1576  XOR n_1580;
or1_1259: n_1576 <=  n_1577;
and2_1260: n_1577 <=  n_1578  AND n_1579;
inv_1261: n_1578  <= TRANSPORT NOT nRD  ;
inv_1262: n_1579  <= TRANSPORT NOT nCS  ;
and1_1263: n_1580 <=  gnd;
dff_1264: DFF_a8251
    PORT MAP ( D => a_N1810_aD, CLK => a_N1810_aCLK, CLRN => a_N1810_aCLRN,
          PRN => vcc, Q => a_N1810_aQ);
delay_1265: a_N1810_aCLRN  <= TRANSPORT nRESET  ;
xor2_1266: a_N1810_aD <=  n_1588  XOR n_1593;
or1_1267: n_1588 <=  n_1589;
and3_1268: n_1589 <=  n_1590  AND n_1591  AND n_1592;
inv_1269: n_1590  <= TRANSPORT NOT a_LC5_C13_aOUT  ;
inv_1270: n_1591  <= TRANSPORT NOT CnD  ;
delay_1271: n_1592  <= TRANSPORT a_SNEN_aNOT_aOUT  ;
and1_1272: n_1593 <=  gnd;
delay_1273: n_1594  <= TRANSPORT nRXC  ;
filter_1274: FILTER_a8251
    PORT MAP (IN1 => n_1594, Y => a_N1810_aCLK);
dff_1275: DFF_a8251
    PORT MAP ( D => a_N1809_aD, CLK => a_N1809_aCLK, CLRN => a_N1809_aCLRN,
          PRN => vcc, Q => a_N1809_aQ);
delay_1276: a_N1809_aCLRN  <= TRANSPORT nRESET  ;
xor2_1277: a_N1809_aD <=  n_1603  XOR n_1606;
or1_1278: n_1603 <=  n_1604;
and1_1279: n_1604 <=  n_1605;
delay_1280: n_1605  <= TRANSPORT a_N1810_aQ  ;
and1_1281: n_1606 <=  gnd;
delay_1282: n_1607  <= TRANSPORT nRXC  ;
filter_1283: FILTER_a8251
    PORT MAP (IN1 => n_1607, Y => a_N1809_aCLK);
delay_1284: a_N102_aOUT  <= TRANSPORT a_N102_aIN  ;
xor2_1285: a_N102_aIN <=  n_1611  XOR n_1620;
or2_1286: n_1611 <=  n_1612  OR n_1616;
and3_1287: n_1612 <=  n_1613  AND n_1614  AND n_1615;
inv_1288: n_1613  <= TRANSPORT NOT a_N83_aOUT  ;
inv_1289: n_1614  <= TRANSPORT NOT a_N1809_aQ  ;
delay_1290: n_1615  <= TRANSPORT nRESET  ;
and3_1291: n_1616 <=  n_1617  AND n_1618  AND n_1619;
inv_1292: n_1617  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1293: n_1618  <= TRANSPORT a_N1810_aQ  ;
delay_1294: n_1619  <= TRANSPORT nRESET  ;
and1_1295: n_1620 <=  gnd;
dff_1296: DFF_a8251
    PORT MAP ( D => a_N2010_aD, CLK => a_N2010_aCLK, CLRN => a_N2010_aCLRN,
          PRN => vcc, Q => a_N2010_aQ);
delay_1297: a_N2010_aCLRN  <= TRANSPORT nRESET  ;
xor2_1298: a_N2010_aD <=  n_1628  XOR n_1637;
or2_1299: n_1628 <=  n_1629  OR n_1632;
and2_1300: n_1629 <=  n_1630  AND n_1631;
delay_1301: n_1630  <= TRANSPORT a_N102_aOUT  ;
delay_1302: n_1631  <= TRANSPORT a_N2010_aQ  ;
and3_1303: n_1632 <=  n_1633  AND n_1635  AND n_1636;
delay_1304: n_1633  <= TRANSPORT a_N655_aOUT  ;
inv_1305: n_1635  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
delay_1306: n_1636  <= TRANSPORT a_N102_aOUT  ;
and1_1307: n_1637 <=  gnd;
delay_1308: n_1638  <= TRANSPORT nRXC  ;
filter_1309: FILTER_a8251
    PORT MAP (IN1 => n_1638, Y => a_N2010_aCLK);
dff_1310: DFF_a8251
    PORT MAP ( D => a_STXRDY_aNOT_aD, CLK => a_STXRDY_aNOT_aCLK, CLRN => a_STXRDY_aNOT_aCLRN,
          PRN => vcc, Q => a_STXRDY_aNOT_aQ);
delay_1311: a_STXRDY_aNOT_aCLRN  <= TRANSPORT nRESET  ;
xor2_1312: a_STXRDY_aNOT_aD <=  n_1647  XOR n_1657;
or2_1313: n_1647 <=  n_1648  OR n_1653;
and3_1314: n_1648 <=  n_1649  AND n_1650  AND n_1652;
delay_1315: n_1649  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_1316: n_1650  <= TRANSPORT a_N77_aNOT_aOUT  ;
delay_1317: n_1652  <= TRANSPORT a_STXRDY_aNOT_aQ  ;
and2_1318: n_1653 <=  n_1654  AND n_1655;
delay_1319: n_1654  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_1320: n_1655  <= TRANSPORT a_N489_aNOT_aOUT  ;
and1_1321: n_1657 <=  gnd;
inv_1322: n_1658  <= TRANSPORT NOT nTXC  ;
filter_1323: FILTER_a8251
    PORT MAP (IN1 => n_1658, Y => a_STXRDY_aNOT_aCLK);
delay_1324: a_N534_aNOT_aOUT  <= TRANSPORT a_N534_aNOT_aIN  ;
xor2_1325: a_N534_aNOT_aIN <=  n_1662  XOR n_1673;
or3_1326: n_1662 <=  n_1663  OR n_1666  OR n_1669;
and2_1327: n_1663 <=  n_1664  AND n_1665;
delay_1328: n_1664  <= TRANSPORT a_N1107_aOUT  ;
delay_1329: n_1665  <= TRANSPORT a_N414_aQ  ;
and2_1330: n_1666 <=  n_1667  AND n_1668;
delay_1331: n_1667  <= TRANSPORT a_SMODE_OUT_F7_G_aQ  ;
inv_1332: n_1668  <= TRANSPORT NOT a_N414_aQ  ;
and2_1333: n_1669 <=  n_1670  AND n_1672;
delay_1334: n_1670  <= TRANSPORT a_N1136_aNOT_aOUT  ;
inv_1335: n_1672  <= TRANSPORT NOT a_N414_aQ  ;
and1_1336: n_1673 <=  gnd;
delay_1337: a_LC3_B14_aOUT  <= TRANSPORT a_LC3_B14_aIN  ;
xor2_1338: a_LC3_B14_aIN <=  n_1676  XOR n_1686;
or3_1339: n_1676 <=  n_1677  OR n_1680  OR n_1683;
and2_1340: n_1677 <=  n_1678  AND n_1679;
delay_1341: n_1678  <= TRANSPORT a_N534_aNOT_aOUT  ;
delay_1342: n_1679  <= TRANSPORT a_STXEMPTY_aNOT_aQ  ;
and2_1343: n_1680 <=  n_1681  AND n_1682;
delay_1344: n_1681  <= TRANSPORT a_STXRDY_aNOT_aQ  ;
delay_1345: n_1682  <= TRANSPORT a_STXEMPTY_aNOT_aQ  ;
and2_1346: n_1683 <=  n_1684  AND n_1685;
delay_1347: n_1684  <= TRANSPORT a_N1128_aNOT_aOUT  ;
delay_1348: n_1685  <= TRANSPORT a_STXEMPTY_aNOT_aQ  ;
and1_1349: n_1686 <=  gnd;
dff_1350: DFF_a8251
    PORT MAP ( D => a_STXEMPTY_aNOT_aD, CLK => a_STXEMPTY_aNOT_aCLK, CLRN => a_STXEMPTY_aNOT_aCLRN,
          PRN => vcc, Q => a_STXEMPTY_aNOT_aQ);
delay_1351: a_STXEMPTY_aNOT_aCLRN  <= TRANSPORT nRESET  ;
xor2_1352: a_STXEMPTY_aNOT_aD <=  n_1693  XOR n_1701;
or2_1353: n_1693 <=  n_1694  OR n_1698;
and3_1354: n_1694 <=  n_1695  AND n_1696  AND n_1697;
delay_1355: n_1695  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_1356: n_1696  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_1357: n_1697  <= TRANSPORT a_LC3_B14_aOUT  ;
and2_1358: n_1698 <=  n_1699  AND n_1700;
delay_1359: n_1699  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_1360: n_1700  <= TRANSPORT a_N489_aNOT_aOUT  ;
and1_1361: n_1701 <=  gnd;
inv_1362: n_1702  <= TRANSPORT NOT nTXC  ;
filter_1363: FILTER_a8251
    PORT MAP (IN1 => n_1702, Y => a_STXEMPTY_aNOT_aCLK);
dff_1364: DFF_a8251
    PORT MAP ( D => a_SRXRDY_aD, CLK => a_SRXRDY_aCLK, CLRN => a_SRXRDY_aCLRN,
          PRN => vcc, Q => a_SRXRDY_aQ);
delay_1365: a_SRXRDY_aCLRN  <= TRANSPORT nRESET  ;
xor2_1366: a_SRXRDY_aD <=  n_1710  XOR n_1718;
or2_1367: n_1710 <=  n_1711  OR n_1714;
and2_1368: n_1711 <=  n_1712  AND n_1713;
delay_1369: n_1712  <= TRANSPORT a_N102_aOUT  ;
delay_1370: n_1713  <= TRANSPORT a_SRXRDY_aQ  ;
and3_1371: n_1714 <=  n_1715  AND n_1716  AND n_1717;
inv_1372: n_1715  <= TRANSPORT NOT a_N83_aOUT  ;
delay_1373: n_1716  <= TRANSPORT a_N79_aNOT_aOUT  ;
delay_1374: n_1717  <= TRANSPORT a_N102_aOUT  ;
and1_1375: n_1718 <=  gnd;
delay_1376: n_1719  <= TRANSPORT nRXC  ;
filter_1377: FILTER_a8251
    PORT MAP (IN1 => n_1719, Y => a_SRXRDY_aCLK);
dff_1378: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F5_G_aD, CLK => a_SCMND_OUT_F5_G_aCLK, CLRN => a_SCMND_OUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F5_G_aQ);
delay_1379: a_SCMND_OUT_F5_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1380: a_SCMND_OUT_F5_G_aD <=  n_1727  XOR n_1736;
or2_1381: n_1727 <=  n_1728  OR n_1732;
and3_1382: n_1728 <=  n_1729  AND n_1730  AND n_1731;
delay_1383: n_1729  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_1384: n_1730  <= TRANSPORT NOT a_N701_aNOT_aOUT  ;
delay_1385: n_1731  <= TRANSPORT a_SCMND_OUT_F5_G_aQ  ;
and3_1386: n_1732 <=  n_1733  AND n_1734  AND n_1735;
delay_1387: n_1733  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1388: n_1734  <= TRANSPORT a_N701_aNOT_aOUT  ;
delay_1389: n_1735  <= TRANSPORT DIN(5)  ;
and1_1390: n_1736 <=  gnd;
delay_1391: n_1737  <= TRANSPORT CLK  ;
filter_1392: FILTER_a8251
    PORT MAP (IN1 => n_1737, Y => a_SCMND_OUT_F5_G_aCLK);
dff_1393: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F1_G_aD, CLK => a_SCMND_OUT_F1_G_aCLK, CLRN => a_SCMND_OUT_F1_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F1_G_aQ);
delay_1394: a_SCMND_OUT_F1_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_1395: a_SCMND_OUT_F1_G_aD <=  n_1745  XOR n_1754;
or2_1396: n_1745 <=  n_1746  OR n_1750;
and3_1397: n_1746 <=  n_1747  AND n_1748  AND n_1749;
delay_1398: n_1747  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_1399: n_1748  <= TRANSPORT NOT a_N701_aNOT_aOUT  ;
delay_1400: n_1749  <= TRANSPORT a_SCMND_OUT_F1_G_aQ  ;
and3_1401: n_1750 <=  n_1751  AND n_1752  AND n_1753;
delay_1402: n_1751  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_1403: n_1752  <= TRANSPORT a_N701_aNOT_aOUT  ;
delay_1404: n_1753  <= TRANSPORT DIN(1)  ;
and1_1405: n_1754 <=  gnd;
delay_1406: n_1755  <= TRANSPORT CLK  ;
filter_1407: FILTER_a8251
    PORT MAP (IN1 => n_1755, Y => a_SCMND_OUT_F1_G_aCLK);
delay_1408: a_G118_aOUT  <= TRANSPORT a_G118_aIN  ;
xor2_1409: a_G118_aIN <=  n_1758  XOR n_1766;
or2_1410: n_1758 <=  n_1759  OR n_1763;
and3_1411: n_1759 <=  n_1760  AND n_1761  AND n_1762;
delay_1412: n_1760  <= TRANSPORT a_SCMND_OUT_F0_G_aQ  ;
delay_1413: n_1761  <= TRANSPORT CnD  ;
inv_1414: n_1762  <= TRANSPORT NOT a_STXRDY_aNOT_aQ  ;
and2_1415: n_1763 <=  n_1764  AND n_1765;
delay_1416: n_1764  <= TRANSPORT a_SRXREG_F0_G_aQ  ;
inv_1417: n_1765  <= TRANSPORT NOT CnD  ;
and1_1418: n_1766 <=  gnd;
delay_1419: a_G701_aOUT  <= TRANSPORT a_G701_aIN  ;
xor2_1420: a_G701_aIN <=  n_1768  XOR n_1775;
or2_1421: n_1768 <=  n_1769  OR n_1772;
and2_1422: n_1769 <=  n_1770  AND n_1771;
delay_1423: n_1770  <= TRANSPORT CnD  ;
delay_1424: n_1771  <= TRANSPORT a_SRXRDY_aQ  ;
and2_1425: n_1772 <=  n_1773  AND n_1774;
delay_1426: n_1773  <= TRANSPORT a_SRXREG_F1_G_aQ  ;
inv_1427: n_1774  <= TRANSPORT NOT CnD  ;
and1_1428: n_1775 <=  gnd;
delay_1429: a_G705_aOUT  <= TRANSPORT a_G705_aIN  ;
xor2_1430: a_G705_aIN <=  n_1777  XOR n_1784;
or2_1431: n_1777 <=  n_1778  OR n_1781;
and2_1432: n_1778 <=  n_1779  AND n_1780;
delay_1433: n_1779  <= TRANSPORT a_SRXREG_F2_G_aQ  ;
inv_1434: n_1780  <= TRANSPORT NOT CnD  ;
and2_1435: n_1781 <=  n_1782  AND n_1783;
delay_1436: n_1782  <= TRANSPORT CnD  ;
inv_1437: n_1783  <= TRANSPORT NOT a_STXEMPTY_aNOT_aQ  ;
and1_1438: n_1784 <=  gnd;
delay_1439: a_G491_aOUT  <= TRANSPORT a_G491_aIN  ;
xor2_1440: a_G491_aIN <=  n_1786  XOR n_1793;
or2_1441: n_1786 <=  n_1787  OR n_1790;
and2_1442: n_1787 <=  n_1788  AND n_1789;
delay_1443: n_1788  <= TRANSPORT a_SRXREG_F3_G_aQ  ;
inv_1444: n_1789  <= TRANSPORT NOT CnD  ;
and2_1445: n_1790 <=  n_1791  AND n_1792;
delay_1446: n_1791  <= TRANSPORT pe_aQ  ;
delay_1447: n_1792  <= TRANSPORT CnD  ;
and1_1448: n_1793 <=  gnd;
delay_1449: a_G495_aOUT  <= TRANSPORT a_G495_aIN  ;
xor2_1450: a_G495_aIN <=  n_1795  XOR n_1802;
or2_1451: n_1795 <=  n_1796  OR n_1799;
and2_1452: n_1796 <=  n_1797  AND n_1798;
delay_1453: n_1797  <= TRANSPORT a_SRXREG_F4_G_aQ  ;
inv_1454: n_1798  <= TRANSPORT NOT CnD  ;
and2_1455: n_1799 <=  n_1800  AND n_1801;
delay_1456: n_1800  <= TRANSPORT oe_aQ  ;
delay_1457: n_1801  <= TRANSPORT CnD  ;
and1_1458: n_1802 <=  gnd;
delay_1459: a_G483_aOUT  <= TRANSPORT a_G483_aIN  ;
xor2_1460: a_G483_aIN <=  n_1804  XOR n_1811;
or2_1461: n_1804 <=  n_1805  OR n_1808;
and2_1462: n_1805 <=  n_1806  AND n_1807;
delay_1463: n_1806  <= TRANSPORT a_SRXREG_F5_G_aQ  ;
inv_1464: n_1807  <= TRANSPORT NOT CnD  ;
and2_1465: n_1808 <=  n_1809  AND n_1810;
delay_1466: n_1809  <= TRANSPORT fe_aQ  ;
delay_1467: n_1810  <= TRANSPORT CnD  ;
and1_1468: n_1811 <=  gnd;
delay_1469: a_SSYN_BRK_aOUT  <= TRANSPORT a_SSYN_BRK_aIN  ;
xor2_1470: a_SSYN_BRK_aIN <=  n_1813  XOR n_1825;
or3_1471: n_1813 <=  n_1814  OR n_1818  OR n_1821;
and2_1472: n_1814 <=  n_1815  AND n_1817;
inv_1473: n_1815  <= TRANSPORT NOT a_N143_aOUT  ;
delay_1474: n_1817  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and2_1475: n_1818 <=  n_1819  AND n_1820;
inv_1476: n_1819  <= TRANSPORT NOT a_N143_aOUT  ;
delay_1477: n_1820  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and3_1478: n_1821 <=  n_1822  AND n_1823  AND n_1824;
inv_1479: n_1822  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
inv_1480: n_1823  <= TRANSPORT NOT a_SMODE_OUT_F1_G_aQ  ;
delay_1481: n_1824  <= TRANSPORT a_N2010_aQ  ;
and1_1482: n_1825 <=  gnd;
delay_1483: a_G514_aOUT  <= TRANSPORT a_G514_aIN  ;
xor2_1484: a_G514_aIN <=  n_1827  XOR n_1834;
or2_1485: n_1827 <=  n_1828  OR n_1831;
and2_1486: n_1828 <=  n_1829  AND n_1830;
delay_1487: n_1829  <= TRANSPORT CnD  ;
delay_1488: n_1830  <= TRANSPORT a_SSYN_BRK_aOUT  ;
and2_1489: n_1831 <=  n_1832  AND n_1833;
delay_1490: n_1832  <= TRANSPORT a_SRXREG_F6_G_aQ  ;
inv_1491: n_1833  <= TRANSPORT NOT CnD  ;
and1_1492: n_1834 <=  gnd;
delay_1493: a_G708_aOUT  <= TRANSPORT a_G708_aIN  ;
xor2_1494: a_G708_aIN <=  n_1837  XOR n_1844;
or2_1495: n_1837 <=  n_1838  OR n_1841;
and2_1496: n_1838 <=  n_1839  AND n_1840;
delay_1497: n_1839  <= TRANSPORT a_SRXREG_F7_G_aQ  ;
inv_1498: n_1840  <= TRANSPORT NOT CnD  ;
and2_1499: n_1841 <=  n_1842  AND n_1843;
delay_1500: n_1842  <= TRANSPORT CnD  ;
inv_1501: n_1843  <= TRANSPORT NOT nDSR  ;
and1_1502: n_1844 <=  gnd;
delay_1503: a_N435_aOUT  <= TRANSPORT a_N435_aIN  ;
xor2_1504: a_N435_aIN <=  n_1847  XOR n_1857;
or3_1505: n_1847 <=  n_1848  OR n_1851  OR n_1854;
and2_1506: n_1848 <=  n_1849  AND n_1850;
delay_1507: n_1849  <= TRANSPORT a_N411_aQ  ;
inv_1508: n_1850  <= TRANSPORT NOT a_N413_aQ  ;
and2_1509: n_1851 <=  n_1852  AND n_1853;
inv_1510: n_1852  <= TRANSPORT NOT a_N414_aQ  ;
inv_1511: n_1853  <= TRANSPORT NOT a_N413_aQ  ;
and2_1512: n_1854 <=  n_1855  AND n_1856;
delay_1513: n_1855  <= TRANSPORT a_N869_aQ  ;
inv_1514: n_1856  <= TRANSPORT NOT a_N414_aQ  ;
and1_1515: n_1857 <=  gnd;
delay_1516: a_N436_aOUT  <= TRANSPORT a_N436_aIN  ;
xor2_1517: a_N436_aIN <=  n_1860  XOR n_1865;
or1_1518: n_1860 <=  n_1861;
and3_1519: n_1861 <=  n_1862  AND n_1863  AND n_1864;
delay_1520: n_1862  <= TRANSPORT a_N868_aQ  ;
delay_1521: n_1863  <= TRANSPORT a_N414_aQ  ;
delay_1522: n_1864  <= TRANSPORT a_N413_aQ  ;
and1_1523: n_1865 <=  gnd;
delay_1524: a_STXD_aOUT  <= TRANSPORT a_STXD_aIN  ;
xor2_1525: a_STXD_aIN <=  n_1867  XOR n_1876;
or4_1526: n_1867 <=  n_1868  OR n_1870  OR n_1872  OR n_1874;
and1_1527: n_1868 <=  n_1869;
delay_1528: n_1869  <= TRANSPORT a_N435_aOUT  ;
and1_1529: n_1870 <=  n_1871;
delay_1530: n_1871  <= TRANSPORT a_N436_aOUT  ;
and1_1531: n_1872 <=  n_1873;
delay_1532: n_1873  <= TRANSPORT a_SCMND_OUT_F3_G_aQ  ;
and1_1533: n_1874 <=  n_1875;
inv_1534: n_1875  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_1535: n_1876 <=  gnd;
delay_1536: a_N1179_aNOT_aOUT  <= TRANSPORT a_N1179_aNOT_aIN  ;
xor2_1537: a_N1179_aNOT_aIN <=  n_1878  XOR n_1883;
or2_1538: n_1878 <=  n_1879  OR n_1881;
and1_1539: n_1879 <=  n_1880;
inv_1540: n_1880  <= TRANSPORT NOT a_N413_aQ  ;
and1_1541: n_1881 <=  n_1882;
delay_1542: n_1882  <= TRANSPORT a_N414_aQ  ;
and1_1543: n_1883 <=  gnd;
delay_1544: a_N76_aNOT_aOUT  <= TRANSPORT a_N76_aNOT_aIN  ;
xor2_1545: a_N76_aNOT_aIN <=  n_1885  XOR n_1890;
or1_1546: n_1885 <=  n_1886;
and3_1547: n_1886 <=  n_1887  AND n_1888  AND n_1889;
inv_1548: n_1887  <= TRANSPORT NOT a_N411_aQ  ;
inv_1549: n_1888  <= TRANSPORT NOT a_N414_aQ  ;
inv_1550: n_1889  <= TRANSPORT NOT a_N413_aQ  ;
and1_1551: n_1890 <=  gnd;
delay_1552: a_N81_aNOT_aOUT  <= TRANSPORT a_N81_aNOT_aIN  ;
xor2_1553: a_N81_aNOT_aIN <=  n_1892  XOR n_1897;
or2_1554: n_1892 <=  n_1893  OR n_1895;
and1_1555: n_1893 <=  n_1894;
delay_1556: n_1894  <= TRANSPORT a_N1904_aQ  ;
and1_1557: n_1895 <=  n_1896;
inv_1558: n_1896  <= TRANSPORT NOT a_N1903_aQ  ;
and1_1559: n_1897 <=  gnd;
delay_1560: a_LC4_B6_aNOT_aOUT  <= TRANSPORT a_LC4_B6_aNOT_aIN  ;
xor2_1561: a_LC4_B6_aNOT_aIN <=  n_1900  XOR n_1907;
or2_1562: n_1900 <=  n_1901  OR n_1904;
and1_1563: n_1901 <=  n_1902;
inv_1564: n_1902  <= TRANSPORT NOT a_N365_aQ  ;
and1_1565: n_1904 <=  n_1905;
inv_1566: n_1905  <= TRANSPORT NOT a_N364_aQ  ;
and1_1567: n_1907 <=  gnd;
delay_1568: a_LC7_B6_aNOT_aOUT  <= TRANSPORT a_LC7_B6_aNOT_aIN  ;
xor2_1569: a_LC7_B6_aNOT_aIN <=  n_1910  XOR n_1916;
or2_1570: n_1910 <=  n_1911  OR n_1914;
and1_1571: n_1911 <=  n_1912;
inv_1572: n_1912  <= TRANSPORT NOT a_N363_aQ  ;
and1_1573: n_1914 <=  n_1915;
delay_1574: n_1915  <= TRANSPORT a_LC4_B6_aNOT_aOUT  ;
and1_1575: n_1916 <=  gnd;
delay_1576: a_LC3_B1_aNOT_aOUT  <= TRANSPORT a_LC3_B1_aNOT_aIN  ;
xor2_1577: a_LC3_B1_aNOT_aIN <=  n_1919  XOR n_1937;
or5_1578: n_1919 <=  n_1920  OR n_1923  OR n_1927  OR n_1931  OR n_1934;
and1_1579: n_1920 <=  n_1921;
inv_1580: n_1921  <= TRANSPORT NOT a_N362_aQ  ;
and2_1581: n_1923 <=  n_1924  AND n_1926;
delay_1582: n_1924  <= TRANSPORT a_N360_aQ  ;
inv_1583: n_1926  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_1584: n_1927 <=  n_1928  AND n_1930;
delay_1585: n_1928  <= TRANSPORT a_N361_aQ  ;
inv_1586: n_1930  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_1587: n_1931 <=  n_1932  AND n_1933;
inv_1588: n_1932  <= TRANSPORT NOT a_N360_aQ  ;
delay_1589: n_1933  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and2_1590: n_1934 <=  n_1935  AND n_1936;
inv_1591: n_1935  <= TRANSPORT NOT a_N361_aQ  ;
delay_1592: n_1936  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and1_1593: n_1937 <=  gnd;
delay_1594: a_N80_aOUT  <= TRANSPORT a_N80_aIN  ;
xor2_1595: a_N80_aIN <=  n_1939  XOR n_1950;
or3_1596: n_1939 <=  n_1940  OR n_1944  OR n_1947;
and2_1597: n_1940 <=  n_1941  AND n_1943;
delay_1598: n_1941  <= TRANSPORT a_N359_aQ  ;
delay_1599: n_1943  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and2_1600: n_1944 <=  n_1945  AND n_1946;
delay_1601: n_1945  <= TRANSPORT a_LC7_B6_aNOT_aOUT  ;
delay_1602: n_1946  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and2_1603: n_1947 <=  n_1948  AND n_1949;
delay_1604: n_1948  <= TRANSPORT a_LC3_B1_aNOT_aOUT  ;
delay_1605: n_1949  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and1_1606: n_1950 <=  gnd;
delay_1607: a_N1136_aNOT_aOUT  <= TRANSPORT a_N1136_aNOT_aIN  ;
xor2_1608: a_N1136_aNOT_aIN <=  n_1952  XOR n_1959;
or3_1609: n_1952 <=  n_1953  OR n_1955  OR n_1957;
and1_1610: n_1953 <=  n_1954;
delay_1611: n_1954  <= TRANSPORT a_N76_aNOT_aOUT  ;
and1_1612: n_1955 <=  n_1956;
inv_1613: n_1956  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_1614: n_1957 <=  n_1958;
delay_1615: n_1958  <= TRANSPORT a_N80_aOUT  ;
and1_1616: n_1959 <=  gnd;
delay_1617: a_N470_aOUT  <= TRANSPORT a_N470_aIN  ;
xor2_1618: a_N470_aIN <=  n_1961  XOR n_1966;
or2_1619: n_1961 <=  n_1962  OR n_1964;
and1_1620: n_1962 <=  n_1963;
delay_1621: n_1963  <= TRANSPORT a_N1179_aNOT_aOUT  ;
and1_1622: n_1964 <=  n_1965;
delay_1623: n_1965  <= TRANSPORT a_N1136_aNOT_aOUT  ;
and1_1624: n_1966 <=  gnd;
delay_1625: a_LC3_B3_aOUT  <= TRANSPORT a_LC3_B3_aIN  ;
xor2_1626: a_LC3_B3_aIN <=  n_1969  XOR n_1974;
or1_1627: n_1969 <=  n_1970;
and2_1628: n_1970 <=  n_1971  AND n_1972;
delay_1629: n_1971  <= TRANSPORT a_N470_aOUT  ;
delay_1630: n_1972  <= TRANSPORT a_N599_aQ  ;
and1_1631: n_1974 <=  gnd;
delay_1632: a_N311_aOUT  <= TRANSPORT a_N311_aIN  ;
xor2_1633: a_N311_aIN <=  n_1977  XOR n_1985;
or3_1634: n_1977 <=  n_1978  OR n_1980  OR n_1982;
and1_1635: n_1978 <=  n_1979;
inv_1636: n_1979  <= TRANSPORT NOT a_N76_aNOT_aOUT  ;
and1_1637: n_1980 <=  n_1981;
inv_1638: n_1981  <= TRANSPORT NOT a_SCMND_OUT_F0_G_aQ  ;
and1_1639: n_1982 <=  n_1983;
delay_1640: n_1983  <= TRANSPORT nCTS  ;
and1_1641: n_1985 <=  gnd;
delay_1642: a_N1064_aNOT_aOUT  <= TRANSPORT a_N1064_aNOT_aIN  ;
xor2_1643: a_N1064_aNOT_aIN <=  n_1988  XOR n_1995;
or3_1644: n_1988 <=  n_1989  OR n_1991  OR n_1993;
and1_1645: n_1989 <=  n_1990;
delay_1646: n_1990  <= TRANSPORT a_N1136_aNOT_aOUT  ;
and1_1647: n_1991 <=  n_1992;
inv_1648: n_1992  <= TRANSPORT NOT a_N413_aQ  ;
and1_1649: n_1993 <=  n_1994;
inv_1650: n_1994  <= TRANSPORT NOT a_N414_aQ  ;
and1_1651: n_1995 <=  gnd;
delay_1652: a_LC1_B4_aNOT_aOUT  <= TRANSPORT a_LC1_B4_aNOT_aIN  ;
xor2_1653: a_LC1_B4_aNOT_aIN <=  n_1997  XOR n_2012;
or4_1654: n_1997 <=  n_1998  OR n_2002  OR n_2005  OR n_2009;
and2_1655: n_1998 <=  n_1999  AND n_2001;
delay_1656: n_1999  <= TRANSPORT a_N396_aQ  ;
inv_1657: n_2001  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and2_1658: n_2002 <=  n_2003  AND n_2004;
inv_1659: n_2003  <= TRANSPORT NOT a_N396_aQ  ;
delay_1660: n_2004  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and2_1661: n_2005 <=  n_2006  AND n_2008;
delay_1662: n_2006  <= TRANSPORT a_N397_aQ  ;
inv_1663: n_2008  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and2_1664: n_2009 <=  n_2010  AND n_2011;
inv_1665: n_2010  <= TRANSPORT NOT a_N397_aQ  ;
delay_1666: n_2011  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_1667: n_2012 <=  gnd;
delay_1668: a_LC8_B4_aNOT_aOUT  <= TRANSPORT a_LC8_B4_aNOT_aIN  ;
xor2_1669: a_LC8_B4_aNOT_aIN <=  n_2014  XOR n_2023;
or4_1670: n_2014 <=  n_2015  OR n_2017  OR n_2019  OR n_2021;
and1_1671: n_2015 <=  n_2016;
delay_1672: n_2016  <= TRANSPORT a_N80_aOUT  ;
and1_1673: n_2017 <=  n_2018;
inv_1674: n_2018  <= TRANSPORT NOT a_N413_aQ  ;
and1_1675: n_2019 <=  n_2020;
inv_1676: n_2020  <= TRANSPORT NOT a_N394_aQ  ;
and1_1677: n_2021 <=  n_2022;
delay_1678: n_2022  <= TRANSPORT a_LC1_B4_aNOT_aOUT  ;
and1_1679: n_2023 <=  gnd;
delay_1680: a_N1056_aOUT  <= TRANSPORT a_N1056_aIN  ;
xor2_1681: a_N1056_aIN <=  n_2026  XOR n_2033;
or3_1682: n_2026 <=  n_2027  OR n_2029  OR n_2031;
and1_1683: n_2027 <=  n_2028;
delay_1684: n_2028  <= TRANSPORT a_LC8_B4_aNOT_aOUT  ;
and1_1685: n_2029 <=  n_2030;
delay_1686: n_2030  <= TRANSPORT a_N414_aQ  ;
and1_1687: n_2031 <=  n_2032;
inv_1688: n_2032  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_1689: n_2033 <=  gnd;
delay_1690: a_N296_aNOT_aOUT  <= TRANSPORT a_N296_aNOT_aIN  ;
xor2_1691: a_N296_aNOT_aIN <=  n_2035  XOR n_2042;
or2_1692: n_2035 <=  n_2036  OR n_2039;
and2_1693: n_2036 <=  n_2037  AND n_2038;
delay_1694: n_2037  <= TRANSPORT a_N1064_aNOT_aOUT  ;
delay_1695: n_2038  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_1696: n_2039 <=  n_2040  AND n_2041;
delay_1697: n_2040  <= TRANSPORT a_N1064_aNOT_aOUT  ;
delay_1698: n_2041  <= TRANSPORT a_N1056_aOUT  ;
and1_1699: n_2042 <=  gnd;
delay_1700: a_N130_aNOT_aOUT  <= TRANSPORT a_N130_aNOT_aIN  ;
xor2_1701: a_N130_aNOT_aIN <=  n_2044  XOR n_2048;
or1_1702: n_2044 <=  n_2045;
and2_1703: n_2045 <=  n_2046  AND n_2047;
inv_1704: n_2046  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
inv_1705: n_2047  <= TRANSPORT NOT a_SMODE_OUT_F1_G_aQ  ;
and1_1706: n_2048 <=  gnd;
delay_1707: a_LC1_B8_aNOT_aOUT  <= TRANSPORT a_LC1_B8_aNOT_aIN  ;
xor2_1708: a_LC1_B8_aNOT_aIN <=  n_2051  XOR n_2058;
or3_1709: n_2051 <=  n_2052  OR n_2054  OR n_2056;
and1_1710: n_2052 <=  n_2053;
inv_1711: n_2053  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_1712: n_2054 <=  n_2055;
delay_1713: n_2055  <= TRANSPORT a_STXRDY_aNOT_aQ  ;
and1_1714: n_2056 <=  n_2057;
inv_1715: n_2057  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
and1_1716: n_2058 <=  gnd;
delay_1717: a_N1114_aNOT_aOUT  <= TRANSPORT a_N1114_aNOT_aIN  ;
xor2_1718: a_N1114_aNOT_aIN <=  n_2060  XOR n_2066;
or2_1719: n_2060 <=  n_2061  OR n_2064;
and2_1720: n_2061 <=  n_2062  AND n_2063;
delay_1721: n_2062  <= TRANSPORT a_N311_aOUT  ;
delay_1722: n_2063  <= TRANSPORT a_N296_aNOT_aOUT  ;
and1_1723: n_2064 <=  n_2065;
delay_1724: n_2065  <= TRANSPORT a_LC1_B8_aNOT_aOUT  ;
and1_1725: n_2066 <=  gnd;
delay_1726: a_LC2_B7_aNOT_aOUT  <= TRANSPORT a_LC2_B7_aNOT_aIN  ;
xor2_1727: a_LC2_B7_aNOT_aIN <=  n_2069  XOR n_2076;
or3_1728: n_2069 <=  n_2070  OR n_2072  OR n_2074;
and1_1729: n_2070 <=  n_2071;
inv_1730: n_2071  <= TRANSPORT NOT a_STXRDY_aNOT_aQ  ;
and1_1731: n_2072 <=  n_2073;
delay_1732: n_2073  <= TRANSPORT a_N413_aQ  ;
and1_1733: n_2074 <=  n_2075;
delay_1734: n_2075  <= TRANSPORT a_N411_aQ  ;
and1_1735: n_2076 <=  gnd;
delay_1736: a_LC3_B7_aNOT_aOUT  <= TRANSPORT a_LC3_B7_aNOT_aIN  ;
xor2_1737: a_LC3_B7_aNOT_aIN <=  n_2078  XOR n_2087;
or4_1738: n_2078 <=  n_2079  OR n_2081  OR n_2083  OR n_2085;
and1_1739: n_2079 <=  n_2080;
inv_1740: n_2080  <= TRANSPORT NOT a_SCMND_OUT_F0_G_aQ  ;
and1_1741: n_2081 <=  n_2082;
delay_1742: n_2082  <= TRANSPORT nCTS  ;
and1_1743: n_2083 <=  n_2084;
delay_1744: n_2084  <= TRANSPORT a_LC2_B7_aNOT_aOUT  ;
and1_1745: n_2085 <=  n_2086;
delay_1746: n_2086  <= TRANSPORT a_N130_aNOT_aOUT  ;
and1_1747: n_2087 <=  gnd;
delay_1748: a_N284_aOUT  <= TRANSPORT a_N284_aIN  ;
xor2_1749: a_N284_aIN <=  n_2090  XOR n_2095;
or2_1750: n_2090 <=  n_2091  OR n_2093;
and1_1751: n_2091 <=  n_2092;
delay_1752: n_2092  <= TRANSPORT a_N414_aQ  ;
and1_1753: n_2093 <=  n_2094;
delay_1754: n_2094  <= TRANSPORT a_LC3_B7_aNOT_aOUT  ;
and1_1755: n_2095 <=  gnd;
delay_1756: a_N1066_aNOT_aOUT  <= TRANSPORT a_N1066_aNOT_aIN  ;
xor2_1757: a_N1066_aNOT_aIN <=  n_2097  XOR n_2104;
or3_1758: n_2097 <=  n_2098  OR n_2100  OR n_2102;
and1_1759: n_2098 <=  n_2099;
inv_1760: n_2099  <= TRANSPORT NOT a_SCMND_OUT_F0_G_aQ  ;
and1_1761: n_2100 <=  n_2101;
delay_1762: n_2101  <= TRANSPORT nCTS  ;
and1_1763: n_2102 <=  n_2103;
inv_1764: n_2103  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
and1_1765: n_2104 <=  gnd;
delay_1766: a_N298_aOUT  <= TRANSPORT a_N298_aIN  ;
xor2_1767: a_N298_aIN <=  n_2106  XOR n_2111;
or2_1768: n_2106 <=  n_2107  OR n_2109;
and1_1769: n_2107 <=  n_2108;
delay_1770: n_2108  <= TRANSPORT a_SMODE_OUT_F7_G_aQ  ;
and1_1771: n_2109 <=  n_2110;
delay_1772: n_2110  <= TRANSPORT a_N80_aOUT  ;
and1_1773: n_2111 <=  gnd;
delay_1774: a_LC2_B16_aNOT_aOUT  <= TRANSPORT a_LC2_B16_aNOT_aIN  ;
xor2_1775: a_LC2_B16_aNOT_aIN <=  n_2114  XOR n_2121;
or3_1776: n_2114 <=  n_2115  OR n_2117  OR n_2119;
and1_1777: n_2115 <=  n_2116;
delay_1778: n_2116  <= TRANSPORT a_N414_aQ  ;
and1_1779: n_2117 <=  n_2118;
delay_1780: n_2118  <= TRANSPORT a_N413_aQ  ;
and1_1781: n_2119 <=  n_2120;
inv_1782: n_2120  <= TRANSPORT NOT a_N411_aQ  ;
and1_1783: n_2121 <=  gnd;
delay_1784: a_LC5_B16_aNOT_aOUT  <= TRANSPORT a_LC5_B16_aNOT_aIN  ;
xor2_1785: a_LC5_B16_aNOT_aIN <=  n_2124  XOR n_2137;
or4_1786: n_2124 <=  n_2125  OR n_2128  OR n_2131  OR n_2134;
and2_1787: n_2125 <=  n_2126  AND n_2127;
delay_1788: n_2126  <= TRANSPORT a_N1066_aNOT_aOUT  ;
delay_1789: n_2127  <= TRANSPORT a_N298_aOUT  ;
and2_1790: n_2128 <=  n_2129  AND n_2130;
delay_1791: n_2129  <= TRANSPORT a_N1066_aNOT_aOUT  ;
delay_1792: n_2130  <= TRANSPORT a_LC2_B16_aNOT_aOUT  ;
and2_1793: n_2131 <=  n_2132  AND n_2133;
inv_1794: n_2132  <= TRANSPORT NOT a_N76_aNOT_aOUT  ;
delay_1795: n_2133  <= TRANSPORT a_N298_aOUT  ;
and2_1796: n_2134 <=  n_2135  AND n_2136;
inv_1797: n_2135  <= TRANSPORT NOT a_N76_aNOT_aOUT  ;
delay_1798: n_2136  <= TRANSPORT a_LC2_B16_aNOT_aOUT  ;
and1_1799: n_2137 <=  gnd;
delay_1800: a_LC6_B1_aNOT_aOUT  <= TRANSPORT a_LC6_B1_aNOT_aIN  ;
xor2_1801: a_LC6_B1_aNOT_aIN <=  n_2140  XOR n_2155;
or5_1802: n_2140 <=  n_2141  OR n_2143  OR n_2146  OR n_2149  OR n_2152;
and1_1803: n_2141 <=  n_2142;
delay_1804: n_2142  <= TRANSPORT a_N360_aQ  ;
and2_1805: n_2143 <=  n_2144  AND n_2145;
delay_1806: n_2144  <= TRANSPORT a_N362_aQ  ;
inv_1807: n_2145  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_1808: n_2146 <=  n_2147  AND n_2148;
delay_1809: n_2147  <= TRANSPORT a_N361_aQ  ;
inv_1810: n_2148  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_1811: n_2149 <=  n_2150  AND n_2151;
inv_1812: n_2150  <= TRANSPORT NOT a_N362_aQ  ;
delay_1813: n_2151  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and2_1814: n_2152 <=  n_2153  AND n_2154;
inv_1815: n_2153  <= TRANSPORT NOT a_N361_aQ  ;
delay_1816: n_2154  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and1_1817: n_2155 <=  gnd;
delay_1818: a_LC4_B17_aNOT_aOUT  <= TRANSPORT a_LC4_B17_aNOT_aIN  ;
xor2_1819: a_LC4_B17_aNOT_aIN <=  n_2158  XOR n_2168;
or3_1820: n_2158 <=  n_2159  OR n_2162  OR n_2165;
and2_1821: n_2159 <=  n_2160  AND n_2161;
delay_1822: n_2160  <= TRANSPORT a_N359_aQ  ;
delay_1823: n_2161  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and2_1824: n_2162 <=  n_2163  AND n_2164;
delay_1825: n_2163  <= TRANSPORT a_LC7_B6_aNOT_aOUT  ;
delay_1826: n_2164  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and2_1827: n_2165 <=  n_2166  AND n_2167;
delay_1828: n_2166  <= TRANSPORT a_LC6_B1_aNOT_aOUT  ;
delay_1829: n_2167  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and1_1830: n_2168 <=  gnd;
delay_1831: a_N1184_aNOT_aOUT  <= TRANSPORT a_N1184_aNOT_aIN  ;
xor2_1832: a_N1184_aNOT_aIN <=  n_2171  XOR n_2176;
or2_1833: n_2171 <=  n_2172  OR n_2174;
and1_1834: n_2172 <=  n_2173;
delay_1835: n_2173  <= TRANSPORT a_N76_aNOT_aOUT  ;
and1_1836: n_2174 <=  n_2175;
inv_1837: n_2175  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_1838: n_2176 <=  gnd;
delay_1839: a_N1107_aOUT  <= TRANSPORT a_N1107_aIN  ;
xor2_1840: a_N1107_aIN <=  n_2178  XOR n_2187;
or3_1841: n_2178 <=  n_2179  OR n_2182  OR n_2185;
and2_1842: n_2179 <=  n_2180  AND n_2181;
delay_1843: n_2180  <= TRANSPORT a_N80_aOUT  ;
delay_1844: n_2181  <= TRANSPORT a_SMODE_OUT_F6_G_aQ  ;
and2_1845: n_2182 <=  n_2183  AND n_2184;
delay_1846: n_2183  <= TRANSPORT a_LC4_B17_aNOT_aOUT  ;
inv_1847: n_2184  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_1848: n_2185 <=  n_2186;
delay_1849: n_2186  <= TRANSPORT a_N1184_aNOT_aOUT  ;
and1_1850: n_2187 <=  gnd;
delay_1851: a_N1128_aNOT_aOUT  <= TRANSPORT a_N1128_aNOT_aIN  ;
xor2_1852: a_N1128_aNOT_aIN <=  n_2189  XOR n_2194;
or2_1853: n_2189 <=  n_2190  OR n_2192;
and1_1854: n_2190 <=  n_2191;
delay_1855: n_2191  <= TRANSPORT a_N413_aQ  ;
and1_1856: n_2192 <=  n_2193;
inv_1857: n_2193  <= TRANSPORT NOT a_N411_aQ  ;
and1_1858: n_2194 <=  gnd;
delay_1859: a_N1065_aOUT  <= TRANSPORT a_N1065_aIN  ;
xor2_1860: a_N1065_aIN <=  n_2197  XOR n_2204;
or3_1861: n_2197 <=  n_2198  OR n_2200  OR n_2202;
and1_1862: n_2198 <=  n_2199;
delay_1863: n_2199  <= TRANSPORT a_N1107_aOUT  ;
and1_1864: n_2200 <=  n_2201;
inv_1865: n_2201  <= TRANSPORT NOT a_N414_aQ  ;
and1_1866: n_2202 <=  n_2203;
delay_1867: n_2203  <= TRANSPORT a_N1128_aNOT_aOUT  ;
and1_1868: n_2204 <=  gnd;
delay_1869: a_LC6_B16_aOUT  <= TRANSPORT a_LC6_B16_aIN  ;
xor2_1870: a_LC6_B16_aIN <=  n_2207  XOR n_2216;
or2_1871: n_2207 <=  n_2208  OR n_2212;
and3_1872: n_2208 <=  n_2209  AND n_2210  AND n_2211;
delay_1873: n_2209  <= TRANSPORT a_N296_aNOT_aOUT  ;
delay_1874: n_2210  <= TRANSPORT a_LC5_B16_aNOT_aOUT  ;
delay_1875: n_2211  <= TRANSPORT a_N1065_aOUT  ;
and3_1876: n_2212 <=  n_2213  AND n_2214  AND n_2215;
inv_1877: n_2213  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_1878: n_2214  <= TRANSPORT a_LC5_B16_aNOT_aOUT  ;
delay_1879: n_2215  <= TRANSPORT a_N1065_aOUT  ;
and1_1880: n_2216 <=  gnd;
delay_1881: a_N77_aNOT_aOUT  <= TRANSPORT a_N77_aNOT_aIN  ;
xor2_1882: a_N77_aNOT_aIN <=  n_2218  XOR n_2225;
or2_1883: n_2218 <=  n_2219  OR n_2222;
and2_1884: n_2219 <=  n_2220  AND n_2221;
delay_1885: n_2220  <= TRANSPORT a_N284_aOUT  ;
inv_1886: n_2221  <= TRANSPORT NOT a_STXRDY_aNOT_aQ  ;
and2_1887: n_2222 <=  n_2223  AND n_2224;
delay_1888: n_2223  <= TRANSPORT a_N284_aOUT  ;
delay_1889: n_2224  <= TRANSPORT a_LC6_B16_aOUT  ;
and1_1890: n_2225 <=  gnd;
delay_1891: a_N1032_aNOT_aOUT  <= TRANSPORT a_N1032_aNOT_aIN  ;
xor2_1892: a_N1032_aNOT_aIN <=  n_2228  XOR n_2233;
or2_1893: n_2228 <=  n_2229  OR n_2231;
and1_1894: n_2229 <=  n_2230;
delay_1895: n_2230  <= TRANSPORT a_N77_aNOT_aOUT  ;
and1_1896: n_2231 <=  n_2232;
inv_1897: n_2232  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_1898: n_2233 <=  gnd;
delay_1899: a_N221_aNOT_aOUT  <= TRANSPORT a_N221_aNOT_aIN  ;
xor2_1900: a_N221_aNOT_aIN <=  n_2235  XOR n_2239;
or1_1901: n_2235 <=  n_2236;
and2_1902: n_2236 <=  n_2237  AND n_2238;
delay_1903: n_2237  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_1904: n_2238  <= TRANSPORT a_N1032_aNOT_aOUT  ;
and1_1905: n_2239 <=  gnd;
delay_1906: a_N1134_aNOT_aOUT  <= TRANSPORT a_N1134_aNOT_aIN  ;
xor2_1907: a_N1134_aNOT_aIN <=  n_2242  XOR n_2247;
or2_1908: n_2242 <=  n_2243  OR n_2245;
and1_1909: n_2243 <=  n_2244;
delay_1910: n_2244  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_1911: n_2245 <=  n_2246;
delay_1912: n_2246  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_1913: n_2247 <=  gnd;
delay_1914: a_LC5_C19_aOUT  <= TRANSPORT a_LC5_C19_aIN  ;
xor2_1915: a_LC5_C19_aIN <=  n_2250  XOR n_2261;
or2_1916: n_2250 <=  n_2251  OR n_2256;
and3_1917: n_2251 <=  n_2252  AND n_2253  AND n_2255;
delay_1918: n_2252  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_1919: n_2253  <= TRANSPORT a_SSYNC1_F7_G_aQ  ;
inv_1920: n_2255  <= TRANSPORT NOT a_N729_aQ  ;
and3_1921: n_2256 <=  n_2257  AND n_2258  AND n_2260;
delay_1922: n_2257  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_1923: n_2258  <= TRANSPORT a_SSYNC2_F7_G_aQ  ;
delay_1924: n_2260  <= TRANSPORT a_N729_aQ  ;
and1_1925: n_2261 <=  gnd;
delay_1926: a_LC4_C19_aOUT  <= TRANSPORT a_LC4_C19_aIN  ;
xor2_1927: a_LC4_C19_aIN <=  n_2264  XOR n_2273;
or2_1928: n_2264 <=  n_2265  OR n_2269;
and3_1929: n_2265 <=  n_2266  AND n_2267  AND n_2268;
delay_1930: n_2266  <= TRANSPORT a_LC5_C19_aOUT  ;
delay_1931: n_2267  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
delay_1932: n_2268  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and3_1933: n_2269 <=  n_2270  AND n_2271  AND n_2272;
delay_1934: n_2270  <= TRANSPORT a_LC5_C19_aOUT  ;
inv_1935: n_2271  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
inv_1936: n_2272  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and1_1937: n_2273 <=  gnd;
delay_1938: a_N1138_aOUT  <= TRANSPORT a_N1138_aIN  ;
xor2_1939: a_N1138_aIN <=  n_2276  XOR n_2280;
or1_1940: n_2276 <=  n_2277;
and2_1941: n_2277 <=  n_2278  AND n_2279;
delay_1942: n_2278  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
delay_1943: n_2279  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_1944: n_2280 <=  gnd;
delay_1945: a_N1108_aNOT_aOUT  <= TRANSPORT a_N1108_aNOT_aIN  ;
xor2_1946: a_N1108_aNOT_aIN <=  n_2282  XOR n_2291;
or2_1947: n_2282 <=  n_2283  OR n_2286;
and2_1948: n_2283 <=  n_2284  AND n_2285;
inv_1949: n_2284  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_1950: n_2285  <= TRANSPORT a_LC4_C19_aOUT  ;
and3_1951: n_2286 <=  n_2287  AND n_2288  AND n_2289;
delay_1952: n_2287  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_1953: n_2288  <= TRANSPORT a_N1138_aOUT  ;
delay_1954: n_2289  <= TRANSPORT a_N2024_aQ  ;
and1_1955: n_2291 <=  gnd;
dff_1956: DFF_a8251
    PORT MAP ( D => a_N599_aD, CLK => a_N599_aCLK, CLRN => a_N599_aCLRN, PRN => vcc,
          Q => a_N599_aQ);
delay_1957: a_N599_aCLRN  <= TRANSPORT nRESET  ;
xor2_1958: a_N599_aD <=  n_2298  XOR n_2307;
or2_1959: n_2298 <=  n_2299  OR n_2303;
and3_1960: n_2299 <=  n_2300  AND n_2301  AND n_2302;
delay_1961: n_2300  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_1962: n_2301  <= TRANSPORT a_LC3_B3_aOUT  ;
delay_1963: n_2302  <= TRANSPORT a_N221_aNOT_aOUT  ;
and3_1964: n_2303 <=  n_2304  AND n_2305  AND n_2306;
delay_1965: n_2304  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_1966: n_2305  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_1967: n_2306  <= TRANSPORT a_N1108_aNOT_aOUT  ;
and1_1968: n_2307 <=  gnd;
inv_1969: n_2308  <= TRANSPORT NOT nTXC  ;
filter_1970: FILTER_a8251
    PORT MAP (IN1 => n_2308, Y => a_N599_aCLK);
delay_1971: a_LC2_B11_aOUT  <= TRANSPORT a_LC2_B11_aIN  ;
xor2_1972: a_LC2_B11_aIN <=  n_2311  XOR n_2315;
or1_1973: n_2311 <=  n_2312;
and2_1974: n_2312 <=  n_2313  AND n_2314;
inv_1975: n_2313  <= TRANSPORT NOT a_N1179_aNOT_aOUT  ;
inv_1976: n_2314  <= TRANSPORT NOT a_N80_aOUT  ;
and1_1977: n_2315 <=  gnd;
delay_1978: a_LC4_B3_aOUT  <= TRANSPORT a_LC4_B3_aIN  ;
xor2_1979: a_LC4_B3_aIN <=  n_2318  XOR n_2326;
or2_1980: n_2318 <=  n_2319  OR n_2323;
and2_1981: n_2319 <=  n_2320  AND n_2321;
delay_1982: n_2320  <= TRANSPORT a_N470_aOUT  ;
delay_1983: n_2321  <= TRANSPORT a_N601_aQ  ;
and2_1984: n_2323 <=  n_2324  AND n_2325;
delay_1985: n_2324  <= TRANSPORT a_N599_aQ  ;
delay_1986: n_2325  <= TRANSPORT a_LC2_B11_aOUT  ;
and1_1987: n_2326 <=  gnd;
delay_1988: a_LC3_C19_aOUT  <= TRANSPORT a_LC3_C19_aIN  ;
xor2_1989: a_LC3_C19_aIN <=  n_2329  XOR n_2338;
or2_1990: n_2329 <=  n_2330  OR n_2334;
and2_1991: n_2330 <=  n_2331  AND n_2333;
delay_1992: n_2331  <= TRANSPORT a_SSYNC2_F6_G_aQ  ;
delay_1993: n_2333  <= TRANSPORT a_N729_aQ  ;
and2_1994: n_2334 <=  n_2335  AND n_2337;
delay_1995: n_2335  <= TRANSPORT a_SSYNC1_F6_G_aQ  ;
inv_1996: n_2337  <= TRANSPORT NOT a_N729_aQ  ;
and1_1997: n_2338 <=  gnd;
delay_1998: a_N1099_aNOT_aOUT  <= TRANSPORT a_N1099_aNOT_aIN  ;
xor2_1999: a_N1099_aNOT_aIN <=  n_2340  XOR n_2350;
or2_2000: n_2340 <=  n_2341  OR n_2346;
and3_2001: n_2341 <=  n_2342  AND n_2343  AND n_2345;
delay_2002: n_2342  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_2003: n_2343  <= TRANSPORT a_N2025_aQ  ;
delay_2004: n_2345  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and3_2005: n_2346 <=  n_2347  AND n_2348  AND n_2349;
inv_2006: n_2347  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_2007: n_2348  <= TRANSPORT a_LC3_C19_aOUT  ;
delay_2008: n_2349  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_2009: n_2350 <=  gnd;
dff_2010: DFF_a8251
    PORT MAP ( D => a_N601_aD, CLK => a_N601_aCLK, CLRN => a_N601_aCLRN, PRN => vcc,
          Q => a_N601_aQ);
delay_2011: a_N601_aCLRN  <= TRANSPORT nRESET  ;
xor2_2012: a_N601_aD <=  n_2357  XOR n_2366;
or2_2013: n_2357 <=  n_2358  OR n_2362;
and3_2014: n_2358 <=  n_2359  AND n_2360  AND n_2361;
delay_2015: n_2359  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_2016: n_2360  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_2017: n_2361  <= TRANSPORT a_LC4_B3_aOUT  ;
and3_2018: n_2362 <=  n_2363  AND n_2364  AND n_2365;
delay_2019: n_2363  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_2020: n_2364  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_2021: n_2365  <= TRANSPORT a_N1099_aNOT_aOUT  ;
and1_2022: n_2366 <=  gnd;
inv_2023: n_2367  <= TRANSPORT NOT nTXC  ;
filter_2024: FILTER_a8251
    PORT MAP (IN1 => n_2367, Y => a_N601_aCLK);
delay_2025: a_LC5_B3_aOUT  <= TRANSPORT a_LC5_B3_aIN  ;
xor2_2026: a_LC5_B3_aIN <=  n_2371  XOR n_2379;
or2_2027: n_2371 <=  n_2372  OR n_2376;
and2_2028: n_2372 <=  n_2373  AND n_2374;
delay_2029: n_2373  <= TRANSPORT a_N470_aOUT  ;
delay_2030: n_2374  <= TRANSPORT a_N602_aQ  ;
and2_2031: n_2376 <=  n_2377  AND n_2378;
delay_2032: n_2377  <= TRANSPORT a_LC2_B11_aOUT  ;
delay_2033: n_2378  <= TRANSPORT a_N601_aQ  ;
and1_2034: n_2379 <=  gnd;
delay_2035: a_N526_aOUT  <= TRANSPORT a_N526_aIN  ;
xor2_2036: a_N526_aIN <=  n_2382  XOR n_2393;
or2_2037: n_2382 <=  n_2383  OR n_2388;
and3_2038: n_2383 <=  n_2384  AND n_2385  AND n_2387;
delay_2039: n_2384  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_2040: n_2385  <= TRANSPORT a_SSYNC1_F5_G_aQ  ;
inv_2041: n_2387  <= TRANSPORT NOT a_N729_aQ  ;
and3_2042: n_2388 <=  n_2389  AND n_2390  AND n_2392;
delay_2043: n_2389  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_2044: n_2390  <= TRANSPORT a_SSYNC2_F5_G_aQ  ;
delay_2045: n_2392  <= TRANSPORT a_N729_aQ  ;
and1_2046: n_2393 <=  gnd;
delay_2047: a_N1098_aNOT_aOUT  <= TRANSPORT a_N1098_aNOT_aIN  ;
xor2_2048: a_N1098_aNOT_aIN <=  n_2395  XOR n_2404;
or2_2049: n_2395 <=  n_2396  OR n_2399;
and2_2050: n_2396 <=  n_2397  AND n_2398;
inv_2051: n_2397  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_2052: n_2398  <= TRANSPORT a_N526_aOUT  ;
and3_2053: n_2399 <=  n_2400  AND n_2401  AND n_2402;
delay_2054: n_2400  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_2055: n_2401  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_2056: n_2402  <= TRANSPORT a_N2026_aQ  ;
and1_2057: n_2404 <=  gnd;
dff_2058: DFF_a8251
    PORT MAP ( D => a_N602_aD, CLK => a_N602_aCLK, CLRN => a_N602_aCLRN, PRN => vcc,
          Q => a_N602_aQ);
delay_2059: a_N602_aCLRN  <= TRANSPORT nRESET  ;
xor2_2060: a_N602_aD <=  n_2411  XOR n_2420;
or2_2061: n_2411 <=  n_2412  OR n_2416;
and3_2062: n_2412 <=  n_2413  AND n_2414  AND n_2415;
delay_2063: n_2413  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_2064: n_2414  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_2065: n_2415  <= TRANSPORT a_LC5_B3_aOUT  ;
and3_2066: n_2416 <=  n_2417  AND n_2418  AND n_2419;
delay_2067: n_2417  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_2068: n_2418  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_2069: n_2419  <= TRANSPORT a_N1098_aNOT_aOUT  ;
and1_2070: n_2420 <=  gnd;
inv_2071: n_2421  <= TRANSPORT NOT nTXC  ;
filter_2072: FILTER_a8251
    PORT MAP (IN1 => n_2421, Y => a_N602_aCLK);
delay_2073: a_LC8_B2_aOUT  <= TRANSPORT a_LC8_B2_aIN  ;
xor2_2074: a_LC8_B2_aIN <=  n_2425  XOR n_2433;
or2_2075: n_2425 <=  n_2426  OR n_2430;
and2_2076: n_2426 <=  n_2427  AND n_2428;
delay_2077: n_2427  <= TRANSPORT a_N470_aOUT  ;
delay_2078: n_2428  <= TRANSPORT a_N603_aQ  ;
and2_2079: n_2430 <=  n_2431  AND n_2432;
delay_2080: n_2431  <= TRANSPORT a_LC2_B11_aOUT  ;
delay_2081: n_2432  <= TRANSPORT a_N602_aQ  ;
and1_2082: n_2433 <=  gnd;
delay_2083: a_LC5_C18_aOUT  <= TRANSPORT a_LC5_C18_aIN  ;
xor2_2084: a_LC5_C18_aIN <=  n_2436  XOR n_2445;
or2_2085: n_2436 <=  n_2437  OR n_2441;
and2_2086: n_2437 <=  n_2438  AND n_2440;
delay_2087: n_2438  <= TRANSPORT a_SSYNC2_F4_G_aQ  ;
delay_2088: n_2440  <= TRANSPORT a_N729_aQ  ;
and2_2089: n_2441 <=  n_2442  AND n_2444;
delay_2090: n_2442  <= TRANSPORT a_SSYNC1_F4_G_aQ  ;
inv_2091: n_2444  <= TRANSPORT NOT a_N729_aQ  ;
and1_2092: n_2445 <=  gnd;
delay_2093: a_N1097_aNOT_aOUT  <= TRANSPORT a_N1097_aNOT_aIN  ;
xor2_2094: a_N1097_aNOT_aIN <=  n_2447  XOR n_2455;
or2_2095: n_2447 <=  n_2448  OR n_2451;
and2_2096: n_2448 <=  n_2449  AND n_2450;
inv_2097: n_2449  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_2098: n_2450  <= TRANSPORT a_LC5_C18_aOUT  ;
and2_2099: n_2451 <=  n_2452  AND n_2453;
delay_2100: n_2452  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_2101: n_2453  <= TRANSPORT a_N2027_aQ  ;
and1_2102: n_2455 <=  gnd;
dff_2103: DFF_a8251
    PORT MAP ( D => a_N603_aD, CLK => a_N603_aCLK, CLRN => a_N603_aCLRN, PRN => vcc,
          Q => a_N603_aQ);
delay_2104: a_N603_aCLRN  <= TRANSPORT nRESET  ;
xor2_2105: a_N603_aD <=  n_2462  XOR n_2471;
or2_2106: n_2462 <=  n_2463  OR n_2467;
and3_2107: n_2463 <=  n_2464  AND n_2465  AND n_2466;
delay_2108: n_2464  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_2109: n_2465  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_2110: n_2466  <= TRANSPORT a_LC8_B2_aOUT  ;
and3_2111: n_2467 <=  n_2468  AND n_2469  AND n_2470;
delay_2112: n_2468  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_2113: n_2469  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_2114: n_2470  <= TRANSPORT a_N1097_aNOT_aOUT  ;
and1_2115: n_2471 <=  gnd;
inv_2116: n_2472  <= TRANSPORT NOT nTXC  ;
filter_2117: FILTER_a8251
    PORT MAP (IN1 => n_2472, Y => a_N603_aCLK);
delay_2118: a_N1175_aNOT_aOUT  <= TRANSPORT a_N1175_aNOT_aIN  ;
xor2_2119: a_N1175_aNOT_aIN <=  n_2476  XOR n_2481;
or2_2120: n_2476 <=  n_2477  OR n_2479;
and1_2121: n_2477 <=  n_2478;
inv_2122: n_2478  <= TRANSPORT NOT a_N64_aQ  ;
and1_2123: n_2479 <=  n_2480;
inv_2124: n_2480  <= TRANSPORT NOT a_N62_aQ  ;
and1_2125: n_2481 <=  gnd;
delay_2126: a_N735_aNOT_aOUT  <= TRANSPORT a_N735_aNOT_aIN  ;
xor2_2127: a_N735_aNOT_aIN <=  n_2484  XOR n_2491;
or3_2128: n_2484 <=  n_2485  OR n_2487  OR n_2489;
and1_2129: n_2485 <=  n_2486;
delay_2130: n_2486  <= TRANSPORT a_N1175_aNOT_aOUT  ;
and1_2131: n_2487 <=  n_2488;
delay_2132: n_2488  <= TRANSPORT a_N63_aQ  ;
and1_2133: n_2489 <=  n_2490;
delay_2134: n_2490  <= TRANSPORT a_N61_aQ  ;
and1_2135: n_2491 <=  gnd;
delay_2136: a_LC5_D17_aOUT  <= TRANSPORT a_LC5_D17_aIN  ;
xor2_2137: a_LC5_D17_aIN <=  n_2494  XOR n_2512;
or5_2138: n_2494 <=  n_2495  OR n_2498  OR n_2502  OR n_2506  OR n_2509;
and1_2139: n_2495 <=  n_2496;
inv_2140: n_2496  <= TRANSPORT NOT a_N30_aQ  ;
and2_2141: n_2498 <=  n_2499  AND n_2501;
delay_2142: n_2499  <= TRANSPORT a_N28_aQ  ;
inv_2143: n_2501  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_2144: n_2502 <=  n_2503  AND n_2504;
delay_2145: n_2503  <= TRANSPORT a_N28_aQ  ;
inv_2146: n_2504  <= TRANSPORT NOT a_N29_aQ  ;
and2_2147: n_2506 <=  n_2507  AND n_2508;
inv_2148: n_2507  <= TRANSPORT NOT a_N28_aQ  ;
delay_2149: n_2508  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and2_2150: n_2509 <=  n_2510  AND n_2511;
inv_2151: n_2510  <= TRANSPORT NOT a_N28_aQ  ;
delay_2152: n_2511  <= TRANSPORT a_N29_aQ  ;
and1_2153: n_2512 <=  gnd;
delay_2154: a_N730_aNOT_aOUT  <= TRANSPORT a_N730_aNOT_aIN  ;
xor2_2155: a_N730_aNOT_aIN <=  n_2515  XOR n_2527;
or4_2156: n_2515 <=  n_2516  OR n_2519  OR n_2522  OR n_2525;
and1_2157: n_2516 <=  n_2517;
inv_2158: n_2517  <= TRANSPORT NOT a_N32_aQ  ;
and1_2159: n_2519 <=  n_2520;
inv_2160: n_2520  <= TRANSPORT NOT a_N31_aQ  ;
and1_2161: n_2522 <=  n_2523;
inv_2162: n_2523  <= TRANSPORT NOT a_N33_aQ  ;
and1_2163: n_2525 <=  n_2526;
delay_2164: n_2526  <= TRANSPORT a_LC5_D17_aOUT  ;
and1_2165: n_2527 <=  gnd;
delay_2166: a_LC2_D14_aOUT  <= TRANSPORT a_LC2_D14_aIN  ;
xor2_2167: a_LC2_D14_aIN <=  n_2530  XOR n_2539;
or4_2168: n_2530 <=  n_2531  OR n_2533  OR n_2535  OR n_2537;
and1_2169: n_2531 <=  n_2532;
inv_2170: n_2532  <= TRANSPORT NOT a_N61_aQ  ;
and1_2171: n_2533 <=  n_2534;
inv_2172: n_2534  <= TRANSPORT NOT a_N64_aQ  ;
and1_2173: n_2535 <=  n_2536;
inv_2174: n_2536  <= TRANSPORT NOT a_N63_aQ  ;
and1_2175: n_2537 <=  n_2538;
delay_2176: n_2538  <= TRANSPORT a_N62_aQ  ;
and1_2177: n_2539 <=  gnd;
delay_2178: a_N83_aOUT  <= TRANSPORT a_N83_aIN  ;
xor2_2179: a_N83_aIN <=  n_2541  XOR n_2545;
or1_2180: n_2541 <=  n_2542;
and2_2181: n_2542 <=  n_2543  AND n_2544;
delay_2182: n_2543  <= TRANSPORT a_N1899_aQ  ;
inv_2183: n_2544  <= TRANSPORT NOT a_N1900_aQ  ;
and1_2184: n_2545 <=  gnd;
delay_2185: a_LC1_D14_aNOT_aOUT  <= TRANSPORT a_LC1_D14_aNOT_aIN  ;
xor2_2186: a_LC1_D14_aNOT_aIN <=  n_2548  XOR n_2558;
or3_2187: n_2548 <=  n_2549  OR n_2552  OR n_2555;
and2_2188: n_2549 <=  n_2550  AND n_2551;
delay_2189: n_2550  <= TRANSPORT a_N735_aNOT_aOUT  ;
delay_2190: n_2551  <= TRANSPORT a_N730_aNOT_aOUT  ;
and2_2191: n_2552 <=  n_2553  AND n_2554;
delay_2192: n_2553  <= TRANSPORT a_N735_aNOT_aOUT  ;
delay_2193: n_2554  <= TRANSPORT a_LC2_D14_aOUT  ;
and2_2194: n_2555 <=  n_2556  AND n_2557;
delay_2195: n_2556  <= TRANSPORT a_N735_aNOT_aOUT  ;
delay_2196: n_2557  <= TRANSPORT a_N83_aOUT  ;
and1_2197: n_2558 <=  gnd;
delay_2198: a_N1118_aNOT_aOUT  <= TRANSPORT a_N1118_aNOT_aIN  ;
xor2_2199: a_N1118_aNOT_aIN <=  n_2561  XOR n_2566;
or2_2200: n_2561 <=  n_2562  OR n_2564;
and1_2201: n_2562 <=  n_2563;
inv_2202: n_2563  <= TRANSPORT NOT a_N63_aQ  ;
and1_2203: n_2564 <=  n_2565;
delay_2204: n_2565  <= TRANSPORT a_N61_aQ  ;
and1_2205: n_2566 <=  gnd;
delay_2206: a_N1149_aNOT_aOUT  <= TRANSPORT a_N1149_aNOT_aIN  ;
xor2_2207: a_N1149_aNOT_aIN <=  n_2569  XOR n_2574;
or2_2208: n_2569 <=  n_2570  OR n_2572;
and1_2209: n_2570 <=  n_2571;
delay_2210: n_2571  <= TRANSPORT a_N61_aQ  ;
and1_2211: n_2572 <=  n_2573;
inv_2212: n_2573  <= TRANSPORT NOT a_N62_aQ  ;
and1_2213: n_2574 <=  gnd;
delay_2214: a_N89_aNOT_aOUT  <= TRANSPORT a_N89_aNOT_aIN  ;
xor2_2215: a_N89_aNOT_aIN <=  n_2577  XOR n_2584;
or3_2216: n_2577 <=  n_2578  OR n_2580  OR n_2582;
and1_2217: n_2578 <=  n_2579;
delay_2218: n_2579  <= TRANSPORT a_N63_aQ  ;
and1_2219: n_2580 <=  n_2581;
delay_2220: n_2581  <= TRANSPORT a_N64_aQ  ;
and1_2221: n_2582 <=  n_2583;
delay_2222: n_2583  <= TRANSPORT a_N1149_aNOT_aOUT  ;
and1_2223: n_2584 <=  gnd;
delay_2224: a_N1163_aNOT_aOUT  <= TRANSPORT a_N1163_aNOT_aIN  ;
xor2_2225: a_N1163_aNOT_aIN <=  n_2586  XOR n_2591;
or2_2226: n_2586 <=  n_2587  OR n_2589;
and1_2227: n_2587 <=  n_2588;
inv_2228: n_2588  <= TRANSPORT NOT a_N63_aQ  ;
and1_2229: n_2589 <=  n_2590;
delay_2230: n_2590  <= TRANSPORT a_N64_aQ  ;
and1_2231: n_2591 <=  gnd;
delay_2232: a_N87_aNOT_aOUT  <= TRANSPORT a_N87_aNOT_aIN  ;
xor2_2233: a_N87_aNOT_aIN <=  n_2594  XOR n_2603;
or4_2234: n_2594 <=  n_2595  OR n_2597  OR n_2599  OR n_2601;
and1_2235: n_2595 <=  n_2596;
delay_2236: n_2596  <= TRANSPORT a_N1163_aNOT_aOUT  ;
and1_2237: n_2597 <=  n_2598;
delay_2238: n_2598  <= TRANSPORT a_N59_aQ  ;
and1_2239: n_2599 <=  n_2600;
delay_2240: n_2600  <= TRANSPORT a_N61_aQ  ;
and1_2241: n_2601 <=  n_2602;
delay_2242: n_2602  <= TRANSPORT a_N62_aQ  ;
and1_2243: n_2603 <=  gnd;
delay_2244: a_N352_aOUT  <= TRANSPORT a_N352_aIN  ;
xor2_2245: a_N352_aIN <=  n_2606  XOR n_2610;
or1_2246: n_2606 <=  n_2607;
and2_2247: n_2607 <=  n_2608  AND n_2609;
delay_2248: n_2608  <= TRANSPORT a_N89_aNOT_aOUT  ;
delay_2249: n_2609  <= TRANSPORT a_N87_aNOT_aOUT  ;
and1_2250: n_2610 <=  gnd;
delay_2251: a_N114_aOUT  <= TRANSPORT a_N114_aIN  ;
xor2_2252: a_N114_aIN <=  n_2613  XOR n_2623;
or3_2253: n_2613 <=  n_2614  OR n_2617  OR n_2620;
and2_2254: n_2614 <=  n_2615  AND n_2616;
delay_2255: n_2615  <= TRANSPORT a_N1118_aNOT_aOUT  ;
delay_2256: n_2616  <= TRANSPORT a_N352_aOUT  ;
and2_2257: n_2617 <=  n_2618  AND n_2619;
delay_2258: n_2618  <= TRANSPORT a_N352_aOUT  ;
inv_2259: n_2619  <= TRANSPORT NOT a_N64_aQ  ;
and2_2260: n_2620 <=  n_2621  AND n_2622;
delay_2261: n_2621  <= TRANSPORT a_N352_aOUT  ;
delay_2262: n_2622  <= TRANSPORT a_N62_aQ  ;
and1_2263: n_2623 <=  gnd;
delay_2264: a_N1144_aNOT_aOUT  <= TRANSPORT a_N1144_aNOT_aIN  ;
xor2_2265: a_N1144_aNOT_aIN <=  n_2626  XOR n_2639;
or4_2266: n_2626 <=  n_2627  OR n_2630  OR n_2633  OR n_2637;
and2_2267: n_2627 <=  n_2628  AND n_2629;
inv_2268: n_2628  <= TRANSPORT NOT a_N61_aQ  ;
inv_2269: n_2629  <= TRANSPORT NOT a_N63_aQ  ;
and2_2270: n_2630 <=  n_2631  AND n_2632;
inv_2271: n_2631  <= TRANSPORT NOT a_N62_aQ  ;
inv_2272: n_2632  <= TRANSPORT NOT a_N61_aQ  ;
and3_2273: n_2633 <=  n_2634  AND n_2635  AND n_2636;
delay_2274: n_2634  <= TRANSPORT a_N62_aQ  ;
delay_2275: n_2635  <= TRANSPORT a_N61_aQ  ;
delay_2276: n_2636  <= TRANSPORT a_N63_aQ  ;
and1_2277: n_2637 <=  n_2638;
delay_2278: n_2638  <= TRANSPORT a_N730_aNOT_aOUT  ;
and1_2279: n_2639 <=  gnd;
delay_2280: a_N95_aNOT_aOUT  <= TRANSPORT a_N95_aNOT_aIN  ;
xor2_2281: a_N95_aNOT_aIN <=  n_2642  XOR n_2647;
or2_2282: n_2642 <=  n_2643  OR n_2645;
and1_2283: n_2643 <=  n_2644;
delay_2284: n_2644  <= TRANSPORT a_N1144_aNOT_aOUT  ;
and1_2285: n_2645 <=  n_2646;
delay_2286: n_2646  <= TRANSPORT a_N83_aOUT  ;
and1_2287: n_2647 <=  gnd;
delay_2288: a_N155_aOUT  <= TRANSPORT a_N155_aIN  ;
xor2_2289: a_N155_aIN <=  n_2650  XOR n_2659;
or4_2290: n_2650 <=  n_2651  OR n_2653  OR n_2655  OR n_2657;
and1_2291: n_2651 <=  n_2652;
delay_2292: n_2652  <= TRANSPORT a_N95_aNOT_aOUT  ;
and1_2293: n_2653 <=  n_2654;
inv_2294: n_2654  <= TRANSPORT NOT a_N63_aQ  ;
and1_2295: n_2655 <=  n_2656;
inv_2296: n_2656  <= TRANSPORT NOT a_N64_aQ  ;
and1_2297: n_2657 <=  n_2658;
delay_2298: n_2658  <= TRANSPORT a_N1149_aNOT_aOUT  ;
and1_2299: n_2659 <=  gnd;
delay_2300: a_LC2_D19_aOUT  <= TRANSPORT a_LC2_D19_aIN  ;
xor2_2301: a_LC2_D19_aIN <=  n_2662  XOR n_2669;
or3_2302: n_2662 <=  n_2663  OR n_2665  OR n_2667;
and1_2303: n_2663 <=  n_2664;
delay_2304: n_2664  <= TRANSPORT a_N59_aQ  ;
and1_2305: n_2665 <=  n_2666;
delay_2306: n_2666  <= TRANSPORT a_N63_aQ  ;
and1_2307: n_2667 <=  n_2668;
delay_2308: n_2668  <= TRANSPORT a_N62_aQ  ;
and1_2309: n_2669 <=  gnd;
delay_2310: a_LC2_D17_aOUT  <= TRANSPORT a_LC2_D17_aIN  ;
xor2_2311: a_LC2_D17_aIN <=  n_2672  XOR n_2687;
or5_2312: n_2672 <=  n_2673  OR n_2675  OR n_2678  OR n_2681  OR n_2684;
and1_2313: n_2673 <=  n_2674;
delay_2314: n_2674  <= TRANSPORT a_N28_aQ  ;
and2_2315: n_2675 <=  n_2676  AND n_2677;
inv_2316: n_2676  <= TRANSPORT NOT a_N30_aQ  ;
delay_2317: n_2677  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
and2_2318: n_2678 <=  n_2679  AND n_2680;
inv_2319: n_2679  <= TRANSPORT NOT a_N30_aQ  ;
delay_2320: n_2680  <= TRANSPORT a_N29_aQ  ;
and2_2321: n_2681 <=  n_2682  AND n_2683;
delay_2322: n_2682  <= TRANSPORT a_N30_aQ  ;
inv_2323: n_2683  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_2324: n_2684 <=  n_2685  AND n_2686;
delay_2325: n_2685  <= TRANSPORT a_N30_aQ  ;
inv_2326: n_2686  <= TRANSPORT NOT a_N29_aQ  ;
and1_2327: n_2687 <=  gnd;
delay_2328: a_LC5_D1_aOUT  <= TRANSPORT a_LC5_D1_aIN  ;
xor2_2329: a_LC5_D1_aIN <=  n_2690  XOR n_2699;
or4_2330: n_2690 <=  n_2691  OR n_2693  OR n_2695  OR n_2697;
and1_2331: n_2691 <=  n_2692;
delay_2332: n_2692  <= TRANSPORT a_LC2_D17_aOUT  ;
and1_2333: n_2693 <=  n_2694;
inv_2334: n_2694  <= TRANSPORT NOT a_N32_aQ  ;
and1_2335: n_2695 <=  n_2696;
inv_2336: n_2696  <= TRANSPORT NOT a_N31_aQ  ;
and1_2337: n_2697 <=  n_2698;
inv_2338: n_2698  <= TRANSPORT NOT a_N33_aQ  ;
and1_2339: n_2699 <=  gnd;
delay_2340: a_N116_aNOT_aOUT  <= TRANSPORT a_N116_aNOT_aIN  ;
xor2_2341: a_N116_aNOT_aIN <=  n_2702  XOR n_2715;
or4_2342: n_2702 <=  n_2703  OR n_2705  OR n_2708  OR n_2711;
and1_2343: n_2703 <=  n_2704;
delay_2344: n_2704  <= TRANSPORT a_LC5_D1_aOUT  ;
and2_2345: n_2705 <=  n_2706  AND n_2707;
inv_2346: n_2706  <= TRANSPORT NOT a_N61_aQ  ;
inv_2347: n_2707  <= TRANSPORT NOT a_N63_aQ  ;
and2_2348: n_2708 <=  n_2709  AND n_2710;
inv_2349: n_2709  <= TRANSPORT NOT a_N62_aQ  ;
inv_2350: n_2710  <= TRANSPORT NOT a_N61_aQ  ;
and3_2351: n_2711 <=  n_2712  AND n_2713  AND n_2714;
delay_2352: n_2712  <= TRANSPORT a_N62_aQ  ;
delay_2353: n_2713  <= TRANSPORT a_N61_aQ  ;
delay_2354: n_2714  <= TRANSPORT a_N63_aQ  ;
and1_2355: n_2715 <=  gnd;
delay_2356: a_N751_aNOT_aOUT  <= TRANSPORT a_N751_aNOT_aIN  ;
xor2_2357: a_N751_aNOT_aIN <=  n_2718  XOR n_2723;
or2_2358: n_2718 <=  n_2719  OR n_2721;
and1_2359: n_2719 <=  n_2720;
delay_2360: n_2720  <= TRANSPORT a_N116_aNOT_aOUT  ;
and1_2361: n_2721 <=  n_2722;
delay_2362: n_2722  <= TRANSPORT a_N83_aOUT  ;
and1_2363: n_2723 <=  gnd;
delay_2364: a_N1137_aNOT_aOUT  <= TRANSPORT a_N1137_aNOT_aIN  ;
xor2_2365: a_N1137_aNOT_aIN <=  n_2726  XOR n_2731;
or2_2366: n_2726 <=  n_2727  OR n_2729;
and1_2367: n_2727 <=  n_2728;
delay_2368: n_2728  <= TRANSPORT a_N64_aQ  ;
and1_2369: n_2729 <=  n_2730;
inv_2370: n_2730  <= TRANSPORT NOT a_N62_aQ  ;
and1_2371: n_2731 <=  gnd;
delay_2372: a_LC4_D15_aOUT  <= TRANSPORT a_LC4_D15_aIN  ;
xor2_2373: a_LC4_D15_aIN <=  n_2734  XOR n_2743;
or4_2374: n_2734 <=  n_2735  OR n_2737  OR n_2739  OR n_2741;
and1_2375: n_2735 <=  n_2736;
delay_2376: n_2736  <= TRANSPORT a_N751_aNOT_aOUT  ;
and1_2377: n_2737 <=  n_2738;
delay_2378: n_2738  <= TRANSPORT a_N1137_aNOT_aOUT  ;
and1_2379: n_2739 <=  n_2740;
delay_2380: n_2740  <= TRANSPORT RXD  ;
and1_2381: n_2741 <=  n_2742;
inv_2382: n_2742  <= TRANSPORT NOT a_N63_aQ  ;
and1_2383: n_2743 <=  gnd;
delay_2384: a_LC1_D15_aOUT  <= TRANSPORT a_LC1_D15_aIN  ;
xor2_2385: a_LC1_D15_aIN <=  n_2746  XOR n_2752;
or2_2386: n_2746 <=  n_2747  OR n_2749;
and1_2387: n_2747 <=  n_2748;
delay_2388: n_2748  <= TRANSPORT a_N61_aQ  ;
and2_2389: n_2749 <=  n_2750  AND n_2751;
delay_2390: n_2750  <= TRANSPORT a_LC2_D19_aOUT  ;
delay_2391: n_2751  <= TRANSPORT a_LC4_D15_aOUT  ;
and1_2392: n_2752 <=  gnd;
delay_2393: a_LC2_D15_aOUT  <= TRANSPORT a_LC2_D15_aIN  ;
xor2_2394: a_LC2_D15_aIN <=  n_2755  XOR n_2761;
or1_2395: n_2755 <=  n_2756;
and4_2396: n_2756 <=  n_2757  AND n_2758  AND n_2759  AND n_2760;
delay_2397: n_2757  <= TRANSPORT a_LC1_D14_aNOT_aOUT  ;
delay_2398: n_2758  <= TRANSPORT a_N114_aOUT  ;
delay_2399: n_2759  <= TRANSPORT a_N155_aOUT  ;
delay_2400: n_2760  <= TRANSPORT a_LC1_D15_aOUT  ;
and1_2401: n_2761 <=  gnd;
delay_2402: a_N1152_aNOT_aOUT  <= TRANSPORT a_N1152_aNOT_aIN  ;
xor2_2403: a_N1152_aNOT_aIN <=  n_2764  XOR n_2769;
or2_2404: n_2764 <=  n_2765  OR n_2767;
and1_2405: n_2765 <=  n_2766;
inv_2406: n_2766  <= TRANSPORT NOT a_N61_aQ  ;
and1_2407: n_2767 <=  n_2768;
inv_2408: n_2768  <= TRANSPORT NOT a_N64_aQ  ;
and1_2409: n_2769 <=  gnd;
delay_2410: a_LC5_D10_aOUT  <= TRANSPORT a_LC5_D10_aIN  ;
xor2_2411: a_LC5_D10_aIN <=  n_2772  XOR n_2781;
or4_2412: n_2772 <=  n_2773  OR n_2775  OR n_2777  OR n_2779;
and1_2413: n_2773 <=  n_2774;
delay_2414: n_2774  <= TRANSPORT a_N1152_aNOT_aOUT  ;
and1_2415: n_2775 <=  n_2776;
delay_2416: n_2776  <= TRANSPORT a_N63_aQ  ;
and1_2417: n_2777 <=  n_2778;
delay_2418: n_2778  <= TRANSPORT a_N62_aQ  ;
and1_2419: n_2779 <=  n_2780;
delay_2420: n_2780  <= TRANSPORT a_N730_aNOT_aOUT  ;
and1_2421: n_2781 <=  gnd;
delay_2422: a_N1183_aNOT_aOUT  <= TRANSPORT a_N1183_aNOT_aIN  ;
xor2_2423: a_N1183_aNOT_aIN <=  n_2783  XOR n_2788;
or2_2424: n_2783 <=  n_2784  OR n_2786;
and1_2425: n_2784 <=  n_2785;
inv_2426: n_2785  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_2427: n_2786 <=  n_2787;
inv_2428: n_2787  <= TRANSPORT NOT a_SMODE_OUT_F7_G_aQ  ;
and1_2429: n_2788 <=  gnd;
delay_2430: a_N209_aOUT  <= TRANSPORT a_N209_aIN  ;
xor2_2431: a_N209_aIN <=  n_2791  XOR n_2804;
or4_2432: n_2791 <=  n_2792  OR n_2795  OR n_2798  OR n_2802;
and2_2433: n_2792 <=  n_2793  AND n_2794;
inv_2434: n_2793  <= TRANSPORT NOT a_N61_aQ  ;
inv_2435: n_2794  <= TRANSPORT NOT a_N63_aQ  ;
and2_2436: n_2795 <=  n_2796  AND n_2797;
inv_2437: n_2796  <= TRANSPORT NOT a_N62_aQ  ;
inv_2438: n_2797  <= TRANSPORT NOT a_N61_aQ  ;
and3_2439: n_2798 <=  n_2799  AND n_2800  AND n_2801;
delay_2440: n_2799  <= TRANSPORT a_N62_aQ  ;
delay_2441: n_2800  <= TRANSPORT a_N61_aQ  ;
delay_2442: n_2801  <= TRANSPORT a_N63_aQ  ;
and1_2443: n_2802 <=  n_2803;
delay_2444: n_2803  <= TRANSPORT a_N83_aOUT  ;
and1_2445: n_2804 <=  gnd;
delay_2446: a_N207_aOUT  <= TRANSPORT a_N207_aIN  ;
xor2_2447: a_N207_aIN <=  n_2807  XOR n_2812;
or2_2448: n_2807 <=  n_2808  OR n_2810;
and1_2449: n_2808 <=  n_2809;
inv_2450: n_2809  <= TRANSPORT NOT a_N33_aQ  ;
and1_2451: n_2810 <=  n_2811;
delay_2452: n_2811  <= TRANSPORT a_N209_aOUT  ;
and1_2453: n_2812 <=  gnd;
delay_2454: a_N193_aNOT_aOUT  <= TRANSPORT a_N193_aNOT_aIN  ;
xor2_2455: a_N193_aNOT_aIN <=  n_2815  XOR n_2822;
or3_2456: n_2815 <=  n_2816  OR n_2818  OR n_2820;
and1_2457: n_2816 <=  n_2817;
inv_2458: n_2817  <= TRANSPORT NOT a_N31_aQ  ;
and1_2459: n_2818 <=  n_2819;
inv_2460: n_2819  <= TRANSPORT NOT a_N32_aQ  ;
and1_2461: n_2820 <=  n_2821;
delay_2462: n_2821  <= TRANSPORT a_N207_aOUT  ;
and1_2463: n_2822 <=  gnd;
delay_2464: a_N153_aOUT  <= TRANSPORT a_N153_aIN  ;
xor2_2465: a_N153_aIN <=  n_2825  XOR n_2834;
or4_2466: n_2825 <=  n_2826  OR n_2828  OR n_2830  OR n_2832;
and1_2467: n_2826 <=  n_2827;
delay_2468: n_2827  <= TRANSPORT a_SMODE_OUT_F6_G_aQ  ;
and1_2469: n_2828 <=  n_2829;
inv_2470: n_2829  <= TRANSPORT NOT a_SMODE_OUT_F7_G_aQ  ;
and1_2471: n_2830 <=  n_2831;
delay_2472: n_2831  <= TRANSPORT a_N116_aNOT_aOUT  ;
and1_2473: n_2832 <=  n_2833;
delay_2474: n_2833  <= TRANSPORT a_N193_aNOT_aOUT  ;
and1_2475: n_2834 <=  gnd;
delay_2476: a_N247_aNOT_aOUT  <= TRANSPORT a_N247_aNOT_aIN  ;
xor2_2477: a_N247_aNOT_aIN <=  n_2837  XOR n_2844;
or3_2478: n_2837 <=  n_2838  OR n_2840  OR n_2842;
and1_2479: n_2838 <=  n_2839;
delay_2480: n_2839  <= TRANSPORT a_N63_aQ  ;
and1_2481: n_2840 <=  n_2841;
inv_2482: n_2841  <= TRANSPORT NOT a_N62_aQ  ;
and1_2483: n_2842 <=  n_2843;
delay_2484: n_2843  <= TRANSPORT a_N1152_aNOT_aOUT  ;
and1_2485: n_2844 <=  gnd;
delay_2486: a_N743_aNOT_aOUT  <= TRANSPORT a_N743_aNOT_aIN  ;
xor2_2487: a_N743_aNOT_aIN <=  n_2847  XOR n_2856;
or2_2488: n_2847 <=  n_2848  OR n_2852;
and3_2489: n_2848 <=  n_2849  AND n_2850  AND n_2851;
delay_2490: n_2849  <= TRANSPORT a_N1183_aNOT_aOUT  ;
delay_2491: n_2850  <= TRANSPORT a_N153_aOUT  ;
inv_2492: n_2851  <= TRANSPORT NOT a_N247_aNOT_aOUT  ;
and3_2493: n_2852 <=  n_2853  AND n_2854  AND n_2855;
delay_2494: n_2853  <= TRANSPORT a_N95_aNOT_aOUT  ;
delay_2495: n_2854  <= TRANSPORT a_N153_aOUT  ;
inv_2496: n_2855  <= TRANSPORT NOT a_N247_aNOT_aOUT  ;
and1_2497: n_2856 <=  gnd;
delay_2498: a_N125_aOUT  <= TRANSPORT a_N125_aIN  ;
xor2_2499: a_N125_aIN <=  n_2859  XOR n_2872;
or4_2500: n_2859 <=  n_2860  OR n_2863  OR n_2866  OR n_2869;
and2_2501: n_2860 <=  n_2861  AND n_2862;
delay_2502: n_2861  <= TRANSPORT a_LC5_D10_aOUT  ;
delay_2503: n_2862  <= TRANSPORT a_N743_aNOT_aOUT  ;
and2_2504: n_2863 <=  n_2864  AND n_2865;
delay_2505: n_2864  <= TRANSPORT a_LC5_D10_aOUT  ;
delay_2506: n_2865  <= TRANSPORT a_N247_aNOT_aOUT  ;
and2_2507: n_2866 <=  n_2867  AND n_2868;
delay_2508: n_2867  <= TRANSPORT a_N209_aOUT  ;
delay_2509: n_2868  <= TRANSPORT a_N743_aNOT_aOUT  ;
and2_2510: n_2869 <=  n_2870  AND n_2871;
delay_2511: n_2870  <= TRANSPORT a_N209_aOUT  ;
delay_2512: n_2871  <= TRANSPORT a_N247_aNOT_aOUT  ;
and1_2513: n_2872 <=  gnd;
delay_2514: a_N341_aOUT  <= TRANSPORT a_N341_aIN  ;
xor2_2515: a_N341_aIN <=  n_2875  XOR n_2881;
or2_2516: n_2875 <=  n_2876  OR n_2879;
and2_2517: n_2876 <=  n_2877  AND n_2878;
delay_2518: n_2877  <= TRANSPORT a_LC2_D15_aOUT  ;
delay_2519: n_2878  <= TRANSPORT a_N125_aOUT  ;
and1_2520: n_2879 <=  n_2880;
delay_2521: n_2880  <= TRANSPORT a_N83_aOUT  ;
and1_2522: n_2881 <=  gnd;
dff_2523: DFF_a8251
    PORT MAP ( D => a_N30_aD, CLK => a_N30_aCLK, CLRN => a_N30_aCLRN, PRN => vcc,
          Q => a_N30_aQ);
delay_2524: a_N30_aCLRN  <= TRANSPORT nRESET  ;
xor2_2525: a_N30_aD <=  n_2888  XOR n_2897;
or2_2526: n_2888 <=  n_2889  OR n_2893;
and3_2527: n_2889 <=  n_2890  AND n_2891  AND n_2892;
delay_2528: n_2890  <= TRANSPORT a_N193_aNOT_aOUT  ;
delay_2529: n_2891  <= TRANSPORT a_N341_aOUT  ;
delay_2530: n_2892  <= TRANSPORT a_N30_aQ  ;
and3_2531: n_2893 <=  n_2894  AND n_2895  AND n_2896;
inv_2532: n_2894  <= TRANSPORT NOT a_N193_aNOT_aOUT  ;
delay_2533: n_2895  <= TRANSPORT a_N341_aOUT  ;
inv_2534: n_2896  <= TRANSPORT NOT a_N30_aQ  ;
and1_2535: n_2897 <=  gnd;
delay_2536: n_2898  <= TRANSPORT nRXC  ;
filter_2537: FILTER_a8251
    PORT MAP (IN1 => n_2898, Y => a_N30_aCLK);
delay_2538: a_N200_aOUT  <= TRANSPORT a_N200_aIN  ;
xor2_2539: a_N200_aIN <=  n_2902  XOR n_2907;
or2_2540: n_2902 <=  n_2903  OR n_2905;
and1_2541: n_2903 <=  n_2904;
inv_2542: n_2904  <= TRANSPORT NOT a_N30_aQ  ;
and1_2543: n_2905 <=  n_2906;
delay_2544: n_2906  <= TRANSPORT a_N193_aNOT_aOUT  ;
and1_2545: n_2907 <=  gnd;
dff_2546: DFF_a8251
    PORT MAP ( D => a_N28_aD, CLK => a_N28_aCLK, CLRN => a_N28_aCLRN, PRN => vcc,
          Q => a_N28_aQ);
delay_2547: a_N28_aCLRN  <= TRANSPORT nRESET  ;
xor2_2548: a_N28_aD <=  n_2914  XOR n_2928;
or3_2549: n_2914 <=  n_2915  OR n_2919  OR n_2923;
and3_2550: n_2915 <=  n_2916  AND n_2917  AND n_2918;
delay_2551: n_2916  <= TRANSPORT a_N341_aOUT  ;
delay_2552: n_2917  <= TRANSPORT a_N200_aOUT  ;
delay_2553: n_2918  <= TRANSPORT a_N28_aQ  ;
and3_2554: n_2919 <=  n_2920  AND n_2921  AND n_2922;
delay_2555: n_2920  <= TRANSPORT a_N341_aOUT  ;
delay_2556: n_2921  <= TRANSPORT a_N28_aQ  ;
inv_2557: n_2922  <= TRANSPORT NOT a_N29_aQ  ;
and4_2558: n_2923 <=  n_2924  AND n_2925  AND n_2926  AND n_2927;
delay_2559: n_2924  <= TRANSPORT a_N341_aOUT  ;
inv_2560: n_2925  <= TRANSPORT NOT a_N200_aOUT  ;
inv_2561: n_2926  <= TRANSPORT NOT a_N28_aQ  ;
delay_2562: n_2927  <= TRANSPORT a_N29_aQ  ;
and1_2563: n_2928 <=  gnd;
delay_2564: n_2929  <= TRANSPORT nRXC  ;
filter_2565: FILTER_a8251
    PORT MAP (IN1 => n_2929, Y => a_N28_aCLK);
dff_2566: DFF_a8251
    PORT MAP ( D => a_N29_aD, CLK => a_N29_aCLK, CLRN => a_N29_aCLRN, PRN => vcc,
          Q => a_N29_aQ);
delay_2567: a_N29_aCLRN  <= TRANSPORT nRESET  ;
xor2_2568: a_N29_aD <=  n_2937  XOR n_2951;
or3_2569: n_2937 <=  n_2938  OR n_2942  OR n_2946;
and3_2570: n_2938 <=  n_2939  AND n_2940  AND n_2941;
delay_2571: n_2939  <= TRANSPORT a_N341_aOUT  ;
inv_2572: n_2940  <= TRANSPORT NOT a_N30_aQ  ;
delay_2573: n_2941  <= TRANSPORT a_N29_aQ  ;
and3_2574: n_2942 <=  n_2943  AND n_2944  AND n_2945;
delay_2575: n_2943  <= TRANSPORT a_N193_aNOT_aOUT  ;
delay_2576: n_2944  <= TRANSPORT a_N341_aOUT  ;
delay_2577: n_2945  <= TRANSPORT a_N29_aQ  ;
and4_2578: n_2946 <=  n_2947  AND n_2948  AND n_2949  AND n_2950;
inv_2579: n_2947  <= TRANSPORT NOT a_N193_aNOT_aOUT  ;
delay_2580: n_2948  <= TRANSPORT a_N341_aOUT  ;
delay_2581: n_2949  <= TRANSPORT a_N30_aQ  ;
inv_2582: n_2950  <= TRANSPORT NOT a_N29_aQ  ;
and1_2583: n_2951 <=  gnd;
delay_2584: n_2952  <= TRANSPORT nRXC  ;
filter_2585: FILTER_a8251
    PORT MAP (IN1 => n_2952, Y => a_N29_aCLK);
delay_2586: a_LC5_B2_aOUT  <= TRANSPORT a_LC5_B2_aIN  ;
xor2_2587: a_LC5_B2_aIN <=  n_2956  XOR n_2964;
or2_2588: n_2956 <=  n_2957  OR n_2961;
and2_2589: n_2957 <=  n_2958  AND n_2959;
delay_2590: n_2958  <= TRANSPORT a_N470_aOUT  ;
delay_2591: n_2959  <= TRANSPORT a_N604_aQ  ;
and2_2592: n_2961 <=  n_2962  AND n_2963;
delay_2593: n_2962  <= TRANSPORT a_LC2_B11_aOUT  ;
delay_2594: n_2963  <= TRANSPORT a_N603_aQ  ;
and1_2595: n_2964 <=  gnd;
delay_2596: a_LC5_C1_aOUT  <= TRANSPORT a_LC5_C1_aIN  ;
xor2_2597: a_LC5_C1_aIN <=  n_2967  XOR n_2976;
or2_2598: n_2967 <=  n_2968  OR n_2972;
and2_2599: n_2968 <=  n_2969  AND n_2971;
delay_2600: n_2969  <= TRANSPORT a_SSYNC2_F3_G_aQ  ;
delay_2601: n_2971  <= TRANSPORT a_N729_aQ  ;
and2_2602: n_2972 <=  n_2973  AND n_2975;
delay_2603: n_2973  <= TRANSPORT a_SSYNC1_F3_G_aQ  ;
inv_2604: n_2975  <= TRANSPORT NOT a_N729_aQ  ;
and1_2605: n_2976 <=  gnd;
delay_2606: a_N1096_aNOT_aOUT  <= TRANSPORT a_N1096_aNOT_aIN  ;
xor2_2607: a_N1096_aNOT_aIN <=  n_2978  XOR n_2986;
or2_2608: n_2978 <=  n_2979  OR n_2982;
and2_2609: n_2979 <=  n_2980  AND n_2981;
inv_2610: n_2980  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_2611: n_2981  <= TRANSPORT a_LC5_C1_aOUT  ;
and2_2612: n_2982 <=  n_2983  AND n_2984;
delay_2613: n_2983  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_2614: n_2984  <= TRANSPORT a_N2028_aQ  ;
and1_2615: n_2986 <=  gnd;
dff_2616: DFF_a8251
    PORT MAP ( D => a_N604_aD, CLK => a_N604_aCLK, CLRN => a_N604_aCLRN, PRN => vcc,
          Q => a_N604_aQ);
delay_2617: a_N604_aCLRN  <= TRANSPORT nRESET  ;
xor2_2618: a_N604_aD <=  n_2993  XOR n_3002;
or2_2619: n_2993 <=  n_2994  OR n_2998;
and3_2620: n_2994 <=  n_2995  AND n_2996  AND n_2997;
delay_2621: n_2995  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_2622: n_2996  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_2623: n_2997  <= TRANSPORT a_LC5_B2_aOUT  ;
and3_2624: n_2998 <=  n_2999  AND n_3000  AND n_3001;
delay_2625: n_2999  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_2626: n_3000  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_2627: n_3001  <= TRANSPORT a_N1096_aNOT_aOUT  ;
and1_2628: n_3002 <=  gnd;
inv_2629: n_3003  <= TRANSPORT NOT nTXC  ;
filter_2630: FILTER_a8251
    PORT MAP (IN1 => n_3003, Y => a_N604_aCLK);
dff_2631: DFF_a8251
    PORT MAP ( D => a_N32_aD, CLK => a_N32_aCLK, CLRN => a_N32_aCLRN, PRN => vcc,
          Q => a_N32_aQ);
delay_2632: a_N32_aCLRN  <= TRANSPORT nRESET  ;
xor2_2633: a_N32_aD <=  n_3011  XOR n_3020;
or2_2634: n_3011 <=  n_3012  OR n_3016;
and3_2635: n_3012 <=  n_3013  AND n_3014  AND n_3015;
delay_2636: n_3013  <= TRANSPORT a_N207_aOUT  ;
delay_2637: n_3014  <= TRANSPORT a_N341_aOUT  ;
delay_2638: n_3015  <= TRANSPORT a_N32_aQ  ;
and3_2639: n_3016 <=  n_3017  AND n_3018  AND n_3019;
inv_2640: n_3017  <= TRANSPORT NOT a_N207_aOUT  ;
delay_2641: n_3018  <= TRANSPORT a_N341_aOUT  ;
inv_2642: n_3019  <= TRANSPORT NOT a_N32_aQ  ;
and1_2643: n_3020 <=  gnd;
delay_2644: n_3021  <= TRANSPORT nRXC  ;
filter_2645: FILTER_a8251
    PORT MAP (IN1 => n_3021, Y => a_N32_aCLK);
dff_2646: DFF_a8251
    PORT MAP ( D => a_N31_aD, CLK => a_N31_aCLK, CLRN => a_N31_aCLRN, PRN => vcc,
          Q => a_N31_aQ);
delay_2647: a_N31_aCLRN  <= TRANSPORT nRESET  ;
xor2_2648: a_N31_aD <=  n_3029  XOR n_3043;
or3_2649: n_3029 <=  n_3030  OR n_3034  OR n_3038;
and3_2650: n_3030 <=  n_3031  AND n_3032  AND n_3033;
delay_2651: n_3031  <= TRANSPORT a_N341_aOUT  ;
inv_2652: n_3032  <= TRANSPORT NOT a_N32_aQ  ;
delay_2653: n_3033  <= TRANSPORT a_N31_aQ  ;
and3_2654: n_3034 <=  n_3035  AND n_3036  AND n_3037;
delay_2655: n_3035  <= TRANSPORT a_N207_aOUT  ;
delay_2656: n_3036  <= TRANSPORT a_N341_aOUT  ;
delay_2657: n_3037  <= TRANSPORT a_N31_aQ  ;
and4_2658: n_3038 <=  n_3039  AND n_3040  AND n_3041  AND n_3042;
inv_2659: n_3039  <= TRANSPORT NOT a_N207_aOUT  ;
delay_2660: n_3040  <= TRANSPORT a_N341_aOUT  ;
delay_2661: n_3041  <= TRANSPORT a_N32_aQ  ;
inv_2662: n_3042  <= TRANSPORT NOT a_N31_aQ  ;
and1_2663: n_3043 <=  gnd;
delay_2664: n_3044  <= TRANSPORT nRXC  ;
filter_2665: FILTER_a8251
    PORT MAP (IN1 => n_3044, Y => a_N31_aCLK);
dff_2666: DFF_a8251
    PORT MAP ( D => a_N33_aD, CLK => a_N33_aCLK, CLRN => a_N33_aCLRN, PRN => vcc,
          Q => a_N33_aQ);
delay_2667: a_N33_aCLRN  <= TRANSPORT nRESET  ;
xor2_2668: a_N33_aD <=  n_3052  XOR n_3061;
or2_2669: n_3052 <=  n_3053  OR n_3057;
and3_2670: n_3053 <=  n_3054  AND n_3055  AND n_3056;
inv_2671: n_3054  <= TRANSPORT NOT a_N209_aOUT  ;
delay_2672: n_3055  <= TRANSPORT a_N341_aOUT  ;
inv_2673: n_3056  <= TRANSPORT NOT a_N33_aQ  ;
and3_2674: n_3057 <=  n_3058  AND n_3059  AND n_3060;
delay_2675: n_3058  <= TRANSPORT a_N209_aOUT  ;
delay_2676: n_3059  <= TRANSPORT a_N341_aOUT  ;
delay_2677: n_3060  <= TRANSPORT a_N33_aQ  ;
and1_2678: n_3061 <=  gnd;
delay_2679: n_3062  <= TRANSPORT nRXC  ;
filter_2680: FILTER_a8251
    PORT MAP (IN1 => n_3062, Y => a_N33_aCLK);
delay_2681: a_N85_aNOT_aOUT  <= TRANSPORT a_N85_aNOT_aIN  ;
xor2_2682: a_N85_aNOT_aIN <=  n_3066  XOR n_3073;
or3_2683: n_3066 <=  n_3067  OR n_3069  OR n_3071;
and1_2684: n_3067 <=  n_3068;
inv_2685: n_3068  <= TRANSPORT NOT a_N414_aQ  ;
and1_2686: n_3069 <=  n_3070;
delay_2687: n_3070  <= TRANSPORT a_N413_aQ  ;
and1_2688: n_3071 <=  n_3072;
delay_2689: n_3072  <= TRANSPORT a_N411_aQ  ;
and1_2690: n_3073 <=  gnd;
delay_2691: a_LC8_B10_aOUT  <= TRANSPORT a_LC8_B10_aIN  ;
xor2_2692: a_LC8_B10_aIN <=  n_3075  XOR n_3088;
or4_2693: n_3075 <=  n_3076  OR n_3079  OR n_3082  OR n_3085;
and2_2694: n_3076 <=  n_3077  AND n_3078;
delay_2695: n_3077  <= TRANSPORT a_N311_aOUT  ;
delay_2696: n_3078  <= TRANSPORT a_N85_aNOT_aOUT  ;
and2_2697: n_3079 <=  n_3080  AND n_3081;
delay_2698: n_3080  <= TRANSPORT a_N1136_aNOT_aOUT  ;
delay_2699: n_3081  <= TRANSPORT a_N311_aOUT  ;
and2_2700: n_3082 <=  n_3083  AND n_3084;
inv_2701: n_3083  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_2702: n_3084  <= TRANSPORT a_N85_aNOT_aOUT  ;
and2_2703: n_3085 <=  n_3086  AND n_3087;
delay_2704: n_3086  <= TRANSPORT a_N1136_aNOT_aOUT  ;
inv_2705: n_3087  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
and1_2706: n_3088 <=  gnd;
delay_2707: a_N522_aNOT_aOUT  <= TRANSPORT a_N522_aNOT_aIN  ;
xor2_2708: a_N522_aNOT_aIN <=  n_3091  XOR n_3100;
or3_2709: n_3091 <=  n_3092  OR n_3095  OR n_3098;
and2_2710: n_3092 <=  n_3093  AND n_3094;
delay_2711: n_3093  <= TRANSPORT a_N1107_aOUT  ;
delay_2712: n_3094  <= TRANSPORT a_N414_aQ  ;
and2_2713: n_3095 <=  n_3096  AND n_3097;
delay_2714: n_3096  <= TRANSPORT a_N1136_aNOT_aOUT  ;
inv_2715: n_3097  <= TRANSPORT NOT a_N414_aQ  ;
and1_2716: n_3098 <=  n_3099;
delay_2717: n_3099  <= TRANSPORT a_N1128_aNOT_aOUT  ;
and1_2718: n_3100 <=  gnd;
delay_2719: a_LC7_B10_aOUT  <= TRANSPORT a_LC7_B10_aIN  ;
xor2_2720: a_LC7_B10_aIN <=  n_3103  XOR n_3109;
or1_2721: n_3103 <=  n_3104;
and4_2722: n_3104 <=  n_3105  AND n_3106  AND n_3107  AND n_3108;
delay_2723: n_3105  <= TRANSPORT a_N470_aOUT  ;
delay_2724: n_3106  <= TRANSPORT a_N1064_aNOT_aOUT  ;
delay_2725: n_3107  <= TRANSPORT a_N284_aOUT  ;
delay_2726: n_3108  <= TRANSPORT a_N522_aNOT_aOUT  ;
and1_2727: n_3109 <=  gnd;
delay_2728: a_LC4_B10_aOUT  <= TRANSPORT a_LC4_B10_aIN  ;
xor2_2729: a_LC4_B10_aIN <=  n_3112  XOR n_3118;
or1_2730: n_3112 <=  n_3113;
and4_2731: n_3113 <=  n_3114  AND n_3115  AND n_3116  AND n_3117;
inv_2732: n_3114  <= TRANSPORT NOT a_N76_aNOT_aOUT  ;
delay_2733: n_3115  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_2734: n_3116  <= TRANSPORT a_LC8_B10_aOUT  ;
delay_2735: n_3117  <= TRANSPORT a_LC7_B10_aOUT  ;
and1_2736: n_3118 <=  gnd;
delay_2737: a_LC1_B10_aOUT  <= TRANSPORT a_LC1_B10_aIN  ;
xor2_2738: a_LC1_B10_aIN <=  n_3121  XOR n_3128;
or2_2739: n_3121 <=  n_3122  OR n_3126;
and3_2740: n_3122 <=  n_3123  AND n_3124  AND n_3125;
delay_2741: n_3123  <= TRANSPORT a_N76_aNOT_aOUT  ;
delay_2742: n_3124  <= TRANSPORT a_LC8_B10_aOUT  ;
delay_2743: n_3125  <= TRANSPORT a_LC7_B10_aOUT  ;
and1_2744: n_3126 <=  n_3127;
inv_2745: n_3127  <= TRANSPORT NOT a_N81_aNOT_aOUT  ;
and1_2746: n_3128 <=  gnd;
dff_2747: DFF_a8251
    PORT MAP ( D => a_N365_aD, CLK => a_N365_aCLK, CLRN => a_N365_aCLRN, PRN => vcc,
          Q => a_N365_aQ);
delay_2748: a_N365_aCLRN  <= TRANSPORT nRESET  ;
xor2_2749: a_N365_aD <=  n_3135  XOR n_3142;
or2_2750: n_3135 <=  n_3136  OR n_3139;
and2_2751: n_3136 <=  n_3137  AND n_3138;
delay_2752: n_3137  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_2753: n_3138  <= TRANSPORT NOT a_N365_aQ  ;
and2_2754: n_3139 <=  n_3140  AND n_3141;
delay_2755: n_3140  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_2756: n_3141  <= TRANSPORT a_N365_aQ  ;
and1_2757: n_3142 <=  gnd;
inv_2758: n_3143  <= TRANSPORT NOT nTXC  ;
filter_2759: FILTER_a8251
    PORT MAP (IN1 => n_3143, Y => a_N365_aCLK);
dff_2760: DFF_a8251
    PORT MAP ( D => a_N364_aD, CLK => a_N364_aCLK, CLRN => a_N364_aCLRN, PRN => vcc,
          Q => a_N364_aQ);
delay_2761: a_N364_aCLRN  <= TRANSPORT nRESET  ;
xor2_2762: a_N364_aD <=  n_3151  XOR n_3163;
or3_2763: n_3151 <=  n_3152  OR n_3156  OR n_3160;
and3_2764: n_3152 <=  n_3153  AND n_3154  AND n_3155;
delay_2765: n_3153  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_2766: n_3154  <= TRANSPORT NOT a_N365_aQ  ;
delay_2767: n_3155  <= TRANSPORT a_N364_aQ  ;
and3_2768: n_3156 <=  n_3157  AND n_3158  AND n_3159;
delay_2769: n_3157  <= TRANSPORT a_LC4_B10_aOUT  ;
delay_2770: n_3158  <= TRANSPORT a_N365_aQ  ;
inv_2771: n_3159  <= TRANSPORT NOT a_N364_aQ  ;
and2_2772: n_3160 <=  n_3161  AND n_3162;
delay_2773: n_3161  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_2774: n_3162  <= TRANSPORT a_N364_aQ  ;
and1_2775: n_3163 <=  gnd;
inv_2776: n_3164  <= TRANSPORT NOT nTXC  ;
filter_2777: FILTER_a8251
    PORT MAP (IN1 => n_3164, Y => a_N364_aCLK);
delay_2778: a_N1189_aOUT  <= TRANSPORT a_N1189_aIN  ;
xor2_2779: a_N1189_aIN <=  n_3167  XOR n_3171;
or1_2780: n_3167 <=  n_3168;
and2_2781: n_3168 <=  n_3169  AND n_3170;
delay_2782: n_3169  <= TRANSPORT a_N1804_aQ  ;
inv_2783: n_3170  <= TRANSPORT NOT a_N1807_aQ  ;
and1_2784: n_3171 <=  gnd;
delay_2785: a_N82_aNOT_aOUT  <= TRANSPORT a_N82_aNOT_aIN  ;
xor2_2786: a_N82_aNOT_aIN <=  n_3173  XOR n_3178;
or2_2787: n_3173 <=  n_3174  OR n_3176;
and1_2788: n_3174 <=  n_3175;
inv_2789: n_3175  <= TRANSPORT NOT a_SCMND_OUT_F6_G_aQ  ;
and1_2790: n_3176 <=  n_3177;
delay_2791: n_3177  <= TRANSPORT a_N1895_aQ  ;
and1_2792: n_3178 <=  gnd;
delay_2793: a_N124_aOUT  <= TRANSPORT a_N124_aIN  ;
xor2_2794: a_N124_aIN <=  n_3181  XOR n_3185;
or1_2795: n_3181 <=  n_3182;
and2_2796: n_3182 <=  n_3183  AND n_3184;
delay_2797: n_3183  <= TRANSPORT a_N1189_aOUT  ;
delay_2798: n_3184  <= TRANSPORT a_N82_aNOT_aOUT  ;
and1_2799: n_3185 <=  gnd;
delay_2800: a_N1035_aOUT  <= TRANSPORT a_N1035_aIN  ;
xor2_2801: a_N1035_aIN <=  n_3188  XOR n_3193;
or1_2802: n_3188 <=  n_3189;
and3_2803: n_3189 <=  n_3190  AND n_3191  AND n_3192;
delay_2804: n_3190  <= TRANSPORT a_N124_aOUT  ;
inv_2805: n_3191  <= TRANSPORT NOT a_N1757_aQ  ;
delay_2806: n_3192  <= TRANSPORT a_N1756_aQ  ;
and1_2807: n_3193 <=  gnd;
delay_2808: a_LC1_C9_aOUT  <= TRANSPORT a_LC1_C9_aIN  ;
xor2_2809: a_LC1_C9_aIN <=  n_3196  XOR n_3202;
or1_2810: n_3196 <=  n_3197;
and4_2811: n_3197 <=  n_3198  AND n_3199  AND n_3200  AND n_3201;
delay_2812: n_3198  <= TRANSPORT a_N1189_aOUT  ;
inv_2813: n_3199  <= TRANSPORT NOT a_N1757_aQ  ;
delay_2814: n_3200  <= TRANSPORT a_N1756_aQ  ;
delay_2815: n_3201  <= TRANSPORT DIN(5)  ;
and1_2816: n_3202 <=  gnd;
dff_2817: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F5_G_aD, CLK => a_SSYNC1_F5_G_aCLK, CLRN => a_SSYNC1_F5_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F5_G_aQ);
delay_2818: a_SSYNC1_F5_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_2819: a_SSYNC1_F5_G_aD <=  n_3209  XOR n_3217;
or2_2820: n_3209 <=  n_3210  OR n_3214;
and3_2821: n_3210 <=  n_3211  AND n_3212  AND n_3213;
delay_2822: n_3211  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_2823: n_3212  <= TRANSPORT NOT a_N1035_aOUT  ;
delay_2824: n_3213  <= TRANSPORT a_SSYNC1_F5_G_aQ  ;
and2_2825: n_3214 <=  n_3215  AND n_3216;
delay_2826: n_3215  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_2827: n_3216  <= TRANSPORT a_LC1_C9_aOUT  ;
and1_2828: n_3217 <=  gnd;
delay_2829: n_3218  <= TRANSPORT CLK  ;
filter_2830: FILTER_a8251
    PORT MAP (IN1 => n_3218, Y => a_SSYNC1_F5_G_aCLK);
dff_2831: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F7_G_aD, CLK => a_SSYNC1_F7_G_aCLK, CLRN => a_SSYNC1_F7_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F7_G_aQ);
delay_2832: a_SSYNC1_F7_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_2833: a_SSYNC1_F7_G_aD <=  n_3226  XOR n_3236;
or2_2834: n_3226 <=  n_3227  OR n_3232;
and3_2835: n_3227 <=  n_3228  AND n_3229  AND n_3230;
delay_2836: n_3228  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_2837: n_3229  <= TRANSPORT a_N1035_aOUT  ;
delay_2838: n_3230  <= TRANSPORT DIN(7)  ;
and3_2839: n_3232 <=  n_3233  AND n_3234  AND n_3235;
delay_2840: n_3233  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_2841: n_3234  <= TRANSPORT NOT a_N1035_aOUT  ;
delay_2842: n_3235  <= TRANSPORT a_SSYNC1_F7_G_aQ  ;
and1_2843: n_3236 <=  gnd;
delay_2844: n_3237  <= TRANSPORT CLK  ;
filter_2845: FILTER_a8251
    PORT MAP (IN1 => n_3237, Y => a_SSYNC1_F7_G_aCLK);
delay_2846: a_LC2_C9_aOUT  <= TRANSPORT a_LC2_C9_aIN  ;
xor2_2847: a_LC2_C9_aIN <=  n_3241  XOR n_3247;
or1_2848: n_3241 <=  n_3242;
and4_2849: n_3242 <=  n_3243  AND n_3244  AND n_3245  AND n_3246;
delay_2850: n_3243  <= TRANSPORT a_N1189_aOUT  ;
delay_2851: n_3244  <= TRANSPORT DIN(6)  ;
inv_2852: n_3245  <= TRANSPORT NOT a_N1757_aQ  ;
delay_2853: n_3246  <= TRANSPORT a_N1756_aQ  ;
and1_2854: n_3247 <=  gnd;
dff_2855: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F6_G_aD, CLK => a_SSYNC1_F6_G_aCLK, CLRN => a_SSYNC1_F6_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F6_G_aQ);
delay_2856: a_SSYNC1_F6_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_2857: a_SSYNC1_F6_G_aD <=  n_3254  XOR n_3262;
or2_2858: n_3254 <=  n_3255  OR n_3259;
and3_2859: n_3255 <=  n_3256  AND n_3257  AND n_3258;
delay_2860: n_3256  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_2861: n_3257  <= TRANSPORT NOT a_N1035_aOUT  ;
delay_2862: n_3258  <= TRANSPORT a_SSYNC1_F6_G_aQ  ;
and2_2863: n_3259 <=  n_3260  AND n_3261;
delay_2864: n_3260  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_2865: n_3261  <= TRANSPORT a_LC2_C9_aOUT  ;
and1_2866: n_3262 <=  gnd;
delay_2867: n_3263  <= TRANSPORT CLK  ;
filter_2868: FILTER_a8251
    PORT MAP (IN1 => n_3263, Y => a_SSYNC1_F6_G_aCLK);
delay_2869: a_LC4_C9_aOUT  <= TRANSPORT a_LC4_C9_aIN  ;
xor2_2870: a_LC4_C9_aIN <=  n_3267  XOR n_3273;
or1_2871: n_3267 <=  n_3268;
and4_2872: n_3268 <=  n_3269  AND n_3270  AND n_3271  AND n_3272;
delay_2873: n_3269  <= TRANSPORT a_N1189_aOUT  ;
delay_2874: n_3270  <= TRANSPORT DIN(4)  ;
inv_2875: n_3271  <= TRANSPORT NOT a_N1757_aQ  ;
delay_2876: n_3272  <= TRANSPORT a_N1756_aQ  ;
and1_2877: n_3273 <=  gnd;
dff_2878: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F4_G_aD, CLK => a_SSYNC1_F4_G_aCLK, CLRN => a_SSYNC1_F4_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F4_G_aQ);
delay_2879: a_SSYNC1_F4_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_2880: a_SSYNC1_F4_G_aD <=  n_3280  XOR n_3288;
or2_2881: n_3280 <=  n_3281  OR n_3285;
and3_2882: n_3281 <=  n_3282  AND n_3283  AND n_3284;
delay_2883: n_3282  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_2884: n_3283  <= TRANSPORT NOT a_N1035_aOUT  ;
delay_2885: n_3284  <= TRANSPORT a_SSYNC1_F4_G_aQ  ;
and2_2886: n_3285 <=  n_3286  AND n_3287;
delay_2887: n_3286  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_2888: n_3287  <= TRANSPORT a_LC4_C9_aOUT  ;
and1_2889: n_3288 <=  gnd;
delay_2890: n_3289  <= TRANSPORT CLK  ;
filter_2891: FILTER_a8251
    PORT MAP (IN1 => n_3289, Y => a_SSYNC1_F4_G_aCLK);
delay_2892: a_LC6_B18_aOUT  <= TRANSPORT a_LC6_B18_aIN  ;
xor2_2893: a_LC6_B18_aIN <=  n_3293  XOR n_3301;
or2_2894: n_3293 <=  n_3294  OR n_3298;
and2_2895: n_3294 <=  n_3295  AND n_3296;
delay_2896: n_3295  <= TRANSPORT a_N470_aOUT  ;
delay_2897: n_3296  <= TRANSPORT a_N605_aQ  ;
and2_2898: n_3298 <=  n_3299  AND n_3300;
delay_2899: n_3299  <= TRANSPORT a_LC2_B11_aOUT  ;
delay_2900: n_3300  <= TRANSPORT a_N604_aQ  ;
and1_2901: n_3301 <=  gnd;
delay_2902: a_LC6_B19_aOUT  <= TRANSPORT a_LC6_B19_aIN  ;
xor2_2903: a_LC6_B19_aIN <=  n_3304  XOR n_3313;
or2_2904: n_3304 <=  n_3305  OR n_3309;
and2_2905: n_3305 <=  n_3306  AND n_3308;
delay_2906: n_3306  <= TRANSPORT a_SSYNC2_F2_G_aQ  ;
delay_2907: n_3308  <= TRANSPORT a_N729_aQ  ;
and2_2908: n_3309 <=  n_3310  AND n_3312;
delay_2909: n_3310  <= TRANSPORT a_SSYNC1_F2_G_aQ  ;
inv_2910: n_3312  <= TRANSPORT NOT a_N729_aQ  ;
and1_2911: n_3313 <=  gnd;
delay_2912: a_N1095_aNOT_aOUT  <= TRANSPORT a_N1095_aNOT_aIN  ;
xor2_2913: a_N1095_aNOT_aIN <=  n_3315  XOR n_3323;
or2_2914: n_3315 <=  n_3316  OR n_3319;
and2_2915: n_3316 <=  n_3317  AND n_3318;
inv_2916: n_3317  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_2917: n_3318  <= TRANSPORT a_LC6_B19_aOUT  ;
and2_2918: n_3319 <=  n_3320  AND n_3321;
delay_2919: n_3320  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_2920: n_3321  <= TRANSPORT a_N2029_aQ  ;
and1_2921: n_3323 <=  gnd;
dff_2922: DFF_a8251
    PORT MAP ( D => a_N605_aD, CLK => a_N605_aCLK, CLRN => a_N605_aCLRN, PRN => vcc,
          Q => a_N605_aQ);
delay_2923: a_N605_aCLRN  <= TRANSPORT nRESET  ;
xor2_2924: a_N605_aD <=  n_3330  XOR n_3339;
or2_2925: n_3330 <=  n_3331  OR n_3335;
and3_2926: n_3331 <=  n_3332  AND n_3333  AND n_3334;
delay_2927: n_3332  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_2928: n_3333  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_2929: n_3334  <= TRANSPORT a_LC6_B18_aOUT  ;
and3_2930: n_3335 <=  n_3336  AND n_3337  AND n_3338;
delay_2931: n_3336  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_2932: n_3337  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_2933: n_3338  <= TRANSPORT a_N1095_aNOT_aOUT  ;
and1_2934: n_3339 <=  gnd;
inv_2935: n_3340  <= TRANSPORT NOT nTXC  ;
filter_2936: FILTER_a8251
    PORT MAP (IN1 => n_3340, Y => a_N605_aCLK);
delay_2937: a_N129_aNOT_aOUT  <= TRANSPORT a_N129_aNOT_aIN  ;
xor2_2938: a_N129_aNOT_aIN <=  n_3344  XOR n_3360;
or4_2939: n_3344 <=  n_3345  OR n_3350  OR n_3354  OR n_3357;
and3_2940: n_3345 <=  n_3346  AND n_3348  AND n_3349;
inv_2941: n_3346  <= TRANSPORT NOT a_N919_aQ  ;
delay_2942: n_3348  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
delay_2943: n_3349  <= TRANSPORT a_SMODE_OUT_F1_G_aQ  ;
and2_2944: n_3350 <=  n_3351  AND n_3353;
delay_2945: n_3351  <= TRANSPORT a_N917_aQ  ;
inv_2946: n_3353  <= TRANSPORT NOT a_SMODE_OUT_F0_G_aQ  ;
and2_2947: n_3354 <=  n_3355  AND n_3356;
delay_2948: n_3355  <= TRANSPORT a_N917_aQ  ;
inv_2949: n_3356  <= TRANSPORT NOT a_SMODE_OUT_F1_G_aQ  ;
and2_2950: n_3357 <=  n_3358  AND n_3359;
delay_2951: n_3358  <= TRANSPORT a_N919_aQ  ;
inv_2952: n_3359  <= TRANSPORT NOT a_N917_aQ  ;
and1_2953: n_3360 <=  gnd;
delay_2954: a_LC8_A9_aOUT  <= TRANSPORT a_LC8_A9_aIN  ;
xor2_2955: a_LC8_A9_aIN <=  n_3363  XOR n_3376;
or4_2956: n_3363 <=  n_3364  OR n_3367  OR n_3370  OR n_3373;
and1_2957: n_3364 <=  n_3365;
inv_2958: n_3365  <= TRANSPORT NOT a_N920_aQ  ;
and1_2959: n_3367 <=  n_3368;
inv_2960: n_3368  <= TRANSPORT NOT a_N923_aQ  ;
and1_2961: n_3370 <=  n_3371;
inv_2962: n_3371  <= TRANSPORT NOT a_N921_aQ  ;
and1_2963: n_3373 <=  n_3374;
inv_2964: n_3374  <= TRANSPORT NOT a_N922_aQ  ;
and1_2965: n_3376 <=  gnd;
delay_2966: a_N1126_aOUT  <= TRANSPORT a_N1126_aIN  ;
xor2_2967: a_N1126_aIN <=  n_3379  XOR n_3388;
or2_2968: n_3379 <=  n_3380  OR n_3384;
and3_2969: n_3380 <=  n_3381  AND n_3382  AND n_3383;
delay_2970: n_3381  <= TRANSPORT a_N129_aNOT_aOUT  ;
delay_2971: n_3382  <= TRANSPORT RXD  ;
delay_2972: n_3383  <= TRANSPORT nRESET  ;
and3_2973: n_3384 <=  n_3385  AND n_3386  AND n_3387;
delay_2974: n_3385  <= TRANSPORT a_LC8_A9_aOUT  ;
delay_2975: n_3386  <= TRANSPORT RXD  ;
delay_2976: n_3387  <= TRANSPORT nRESET  ;
and1_2977: n_3388 <=  gnd;
dff_2978: DFF_a8251
    PORT MAP ( D => a_N919_aD, CLK => a_N919_aCLK, CLRN => a_N919_aCLRN, PRN => vcc,
          Q => a_N919_aQ);
delay_2979: a_N919_aCLRN  <= TRANSPORT nRESET  ;
xor2_2980: a_N919_aD <=  n_3395  XOR n_3410;
or3_2981: n_3395 <=  n_3396  OR n_3401  OR n_3405;
and3_2982: n_3396 <=  n_3397  AND n_3398  AND n_3399;
delay_2983: n_3397  <= TRANSPORT a_N1126_aOUT  ;
delay_2984: n_3398  <= TRANSPORT a_N919_aQ  ;
inv_2985: n_3399  <= TRANSPORT NOT a_SCMND_OUT_F2_G_aQ  ;
and3_2986: n_3401 <=  n_3402  AND n_3403  AND n_3404;
delay_2987: n_3402  <= TRANSPORT a_LC8_A9_aOUT  ;
delay_2988: n_3403  <= TRANSPORT a_N1126_aOUT  ;
delay_2989: n_3404  <= TRANSPORT a_N919_aQ  ;
and4_2990: n_3405 <=  n_3406  AND n_3407  AND n_3408  AND n_3409;
inv_2991: n_3406  <= TRANSPORT NOT a_LC8_A9_aOUT  ;
delay_2992: n_3407  <= TRANSPORT a_N1126_aOUT  ;
inv_2993: n_3408  <= TRANSPORT NOT a_N919_aQ  ;
delay_2994: n_3409  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_2995: n_3410 <=  gnd;
inv_2996: n_3411  <= TRANSPORT NOT nRXC  ;
filter_2997: FILTER_a8251
    PORT MAP (IN1 => n_3411, Y => a_N919_aCLK);
delay_2998: a_N576_aOUT  <= TRANSPORT a_N576_aIN  ;
xor2_2999: a_N576_aIN <=  n_3415  XOR n_3420;
or1_3000: n_3415 <=  n_3416;
and3_3001: n_3416 <=  n_3417  AND n_3418  AND n_3419;
delay_3002: n_3417  <= TRANSPORT a_N923_aQ  ;
delay_3003: n_3418  <= TRANSPORT a_N922_aQ  ;
delay_3004: n_3419  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_3005: n_3420 <=  gnd;
delay_3006: a_N564_aOUT  <= TRANSPORT a_N564_aIN  ;
xor2_3007: a_N564_aIN <=  n_3423  XOR n_3429;
or1_3008: n_3423 <=  n_3424;
and4_3009: n_3424 <=  n_3425  AND n_3426  AND n_3427  AND n_3428;
delay_3010: n_3425  <= TRANSPORT a_N919_aQ  ;
delay_3011: n_3426  <= TRANSPORT a_N576_aOUT  ;
delay_3012: n_3427  <= TRANSPORT a_N920_aQ  ;
delay_3013: n_3428  <= TRANSPORT a_N921_aQ  ;
and1_3014: n_3429 <=  gnd;
delay_3015: a_N1083_aOUT  <= TRANSPORT a_N1083_aIN  ;
xor2_3016: a_N1083_aIN <=  n_3432  XOR n_3437;
or2_3017: n_3432 <=  n_3433  OR n_3435;
and1_3018: n_3433 <=  n_3434;
delay_3019: n_3434  <= TRANSPORT a_N129_aNOT_aOUT  ;
and1_3020: n_3435 <=  n_3436;
delay_3021: n_3436  <= TRANSPORT a_LC8_A9_aOUT  ;
and1_3022: n_3437 <=  gnd;
dff_3023: DFF_a8251
    PORT MAP ( D => a_N917_aD, CLK => a_N917_aCLK, CLRN => a_N917_aCLRN, PRN => vcc,
          Q => a_N917_aQ);
delay_3024: a_N917_aCLRN  <= TRANSPORT nRESET  ;
xor2_3025: a_N917_aD <=  n_3444  XOR n_3455;
or2_3026: n_3444 <=  n_3445  OR n_3450;
and4_3027: n_3445 <=  n_3446  AND n_3447  AND n_3448  AND n_3449;
inv_3028: n_3446  <= TRANSPORT NOT a_N564_aOUT  ;
delay_3029: n_3447  <= TRANSPORT a_N1083_aOUT  ;
delay_3030: n_3448  <= TRANSPORT a_N917_aQ  ;
delay_3031: n_3449  <= TRANSPORT RXD  ;
and4_3032: n_3450 <=  n_3451  AND n_3452  AND n_3453  AND n_3454;
delay_3033: n_3451  <= TRANSPORT a_N564_aOUT  ;
delay_3034: n_3452  <= TRANSPORT a_N1083_aOUT  ;
inv_3035: n_3453  <= TRANSPORT NOT a_N917_aQ  ;
delay_3036: n_3454  <= TRANSPORT RXD  ;
and1_3037: n_3455 <=  gnd;
inv_3038: n_3456  <= TRANSPORT NOT nRXC  ;
filter_3039: FILTER_a8251
    PORT MAP (IN1 => n_3456, Y => a_N917_aCLK);
delay_3040: a_LC5_A9_aOUT  <= TRANSPORT a_LC5_A9_aIN  ;
xor2_3041: a_LC5_A9_aIN <=  n_3460  XOR n_3465;
or1_3042: n_3460 <=  n_3461;
and3_3043: n_3461 <=  n_3462  AND n_3463  AND n_3464;
delay_3044: n_3462  <= TRANSPORT a_N923_aQ  ;
delay_3045: n_3463  <= TRANSPORT a_N921_aQ  ;
delay_3046: n_3464  <= TRANSPORT a_N922_aQ  ;
and1_3047: n_3465 <=  gnd;
delay_3048: a_LC6_A9_aOUT  <= TRANSPORT a_LC6_A9_aIN  ;
xor2_3049: a_LC6_A9_aIN <=  n_3468  XOR n_3480;
or3_3050: n_3468 <=  n_3469  OR n_3473  OR n_3476;
and3_3051: n_3469 <=  n_3470  AND n_3471  AND n_3472;
delay_3052: n_3470  <= TRANSPORT a_N129_aNOT_aOUT  ;
delay_3053: n_3471  <= TRANSPORT a_N920_aQ  ;
inv_3054: n_3472  <= TRANSPORT NOT a_SCMND_OUT_F2_G_aQ  ;
and2_3055: n_3473 <=  n_3474  AND n_3475;
inv_3056: n_3474  <= TRANSPORT NOT a_LC5_A9_aOUT  ;
delay_3057: n_3475  <= TRANSPORT a_N920_aQ  ;
and3_3058: n_3476 <=  n_3477  AND n_3478  AND n_3479;
delay_3059: n_3477  <= TRANSPORT a_LC5_A9_aOUT  ;
inv_3060: n_3478  <= TRANSPORT NOT a_N920_aQ  ;
delay_3061: n_3479  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_3062: n_3480 <=  gnd;
dff_3063: DFF_a8251
    PORT MAP ( D => a_N920_aD, CLK => a_N920_aCLK, CLRN => a_N920_aCLRN, PRN => vcc,
          Q => a_N920_aQ);
delay_3064: a_N920_aCLRN  <= TRANSPORT nRESET  ;
xor2_3065: a_N920_aD <=  n_3487  XOR n_3491;
or1_3066: n_3487 <=  n_3488;
and2_3067: n_3488 <=  n_3489  AND n_3490;
delay_3068: n_3489  <= TRANSPORT a_LC6_A9_aOUT  ;
delay_3069: n_3490  <= TRANSPORT RXD  ;
and1_3070: n_3491 <=  gnd;
inv_3071: n_3492  <= TRANSPORT NOT nRXC  ;
filter_3072: FILTER_a8251
    PORT MAP (IN1 => n_3492, Y => a_N920_aCLK);
dff_3073: DFF_a8251
    PORT MAP ( D => a_N923_aD, CLK => a_N923_aCLK, CLRN => a_N923_aCLRN, PRN => vcc,
          Q => a_N923_aQ);
delay_3074: a_N923_aCLRN  <= TRANSPORT nRESET  ;
xor2_3075: a_N923_aD <=  n_3500  XOR n_3509;
or2_3076: n_3500 <=  n_3501  OR n_3505;
and3_3077: n_3501 <=  n_3502  AND n_3503  AND n_3504;
delay_3078: n_3502  <= TRANSPORT a_N1126_aOUT  ;
inv_3079: n_3503  <= TRANSPORT NOT a_N923_aQ  ;
delay_3080: n_3504  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and3_3081: n_3505 <=  n_3506  AND n_3507  AND n_3508;
delay_3082: n_3506  <= TRANSPORT a_N1126_aOUT  ;
delay_3083: n_3507  <= TRANSPORT a_N923_aQ  ;
inv_3084: n_3508  <= TRANSPORT NOT a_SCMND_OUT_F2_G_aQ  ;
and1_3085: n_3509 <=  gnd;
inv_3086: n_3510  <= TRANSPORT NOT nRXC  ;
filter_3087: FILTER_a8251
    PORT MAP (IN1 => n_3510, Y => a_N923_aCLK);
dff_3088: DFF_a8251
    PORT MAP ( D => a_N921_aD, CLK => a_N921_aCLK, CLRN => a_N921_aCLRN, PRN => vcc,
          Q => a_N921_aQ);
delay_3089: a_N921_aCLRN  <= TRANSPORT nRESET  ;
xor2_3090: a_N921_aD <=  n_3518  XOR n_3527;
or2_3091: n_3518 <=  n_3519  OR n_3523;
and3_3092: n_3519 <=  n_3520  AND n_3521  AND n_3522;
delay_3093: n_3520  <= TRANSPORT a_N1126_aOUT  ;
inv_3094: n_3521  <= TRANSPORT NOT a_N576_aOUT  ;
delay_3095: n_3522  <= TRANSPORT a_N921_aQ  ;
and3_3096: n_3523 <=  n_3524  AND n_3525  AND n_3526;
delay_3097: n_3524  <= TRANSPORT a_N1126_aOUT  ;
delay_3098: n_3525  <= TRANSPORT a_N576_aOUT  ;
inv_3099: n_3526  <= TRANSPORT NOT a_N921_aQ  ;
and1_3100: n_3527 <=  gnd;
inv_3101: n_3528  <= TRANSPORT NOT nRXC  ;
filter_3102: FILTER_a8251
    PORT MAP (IN1 => n_3528, Y => a_N921_aCLK);
dff_3103: DFF_a8251
    PORT MAP ( D => a_N922_aD, CLK => a_N922_aCLK, CLRN => a_N922_aCLRN, PRN => vcc,
          Q => a_N922_aQ);
delay_3104: a_N922_aCLRN  <= TRANSPORT nRESET  ;
xor2_3105: a_N922_aD <=  n_3536  XOR n_3550;
or3_3106: n_3536 <=  n_3537  OR n_3541  OR n_3545;
and3_3107: n_3537 <=  n_3538  AND n_3539  AND n_3540;
delay_3108: n_3538  <= TRANSPORT a_N1126_aOUT  ;
delay_3109: n_3539  <= TRANSPORT a_N922_aQ  ;
inv_3110: n_3540  <= TRANSPORT NOT a_SCMND_OUT_F2_G_aQ  ;
and3_3111: n_3541 <=  n_3542  AND n_3543  AND n_3544;
delay_3112: n_3542  <= TRANSPORT a_N1126_aOUT  ;
inv_3113: n_3543  <= TRANSPORT NOT a_N923_aQ  ;
delay_3114: n_3544  <= TRANSPORT a_N922_aQ  ;
and4_3115: n_3545 <=  n_3546  AND n_3547  AND n_3548  AND n_3549;
delay_3116: n_3546  <= TRANSPORT a_N1126_aOUT  ;
delay_3117: n_3547  <= TRANSPORT a_N923_aQ  ;
inv_3118: n_3548  <= TRANSPORT NOT a_N922_aQ  ;
delay_3119: n_3549  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_3120: n_3550 <=  gnd;
inv_3121: n_3551  <= TRANSPORT NOT nRXC  ;
filter_3122: FILTER_a8251
    PORT MAP (IN1 => n_3551, Y => a_N922_aCLK);
delay_3123: a_N489_aNOT_aOUT  <= TRANSPORT a_N489_aNOT_aIN  ;
xor2_3124: a_N489_aNOT_aIN <=  n_3554  XOR n_3558;
or1_3125: n_3554 <=  n_3555;
and2_3126: n_3555 <=  n_3556  AND n_3557;
delay_3127: n_3556  <= TRANSPORT a_N1811_aQ  ;
inv_3128: n_3557  <= TRANSPORT NOT a_N1812_aQ  ;
and1_3129: n_3558 <=  gnd;
delay_3130: a_N1197_aOUT  <= TRANSPORT a_N1197_aIN  ;
xor2_3131: a_N1197_aIN <=  n_3561  XOR n_3566;
or1_3132: n_3561 <=  n_3562;
and3_3133: n_3562 <=  n_3563  AND n_3564  AND n_3565;
delay_3134: n_3563  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_3135: n_3564  <= TRANSPORT a_N489_aNOT_aOUT  ;
delay_3136: n_3565  <= TRANSPORT nRESET  ;
and1_3137: n_3566 <=  gnd;
delay_3138: a_N1198_aOUT  <= TRANSPORT a_N1198_aIN  ;
xor2_3139: a_N1198_aIN <=  n_3569  XOR n_3574;
or1_3140: n_3569 <=  n_3570;
and3_3141: n_3570 <=  n_3571  AND n_3572  AND n_3573;
delay_3142: n_3571  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_3143: n_3572  <= TRANSPORT NOT a_N489_aNOT_aOUT  ;
delay_3144: n_3573  <= TRANSPORT nRESET  ;
and1_3145: n_3574 <=  gnd;
dff_3146: DFF_a8251
    PORT MAP ( D => a_N2027_aD, CLK => a_N2027_aCLK, CLRN => a_N2027_aCLRN,
          PRN => vcc, Q => a_N2027_aQ);
delay_3147: a_N2027_aCLRN  <= TRANSPORT nRESET  ;
xor2_3148: a_N2027_aD <=  n_3581  XOR n_3588;
or2_3149: n_3581 <=  n_3582  OR n_3585;
and2_3150: n_3582 <=  n_3583  AND n_3584;
delay_3151: n_3583  <= TRANSPORT a_N1197_aOUT  ;
delay_3152: n_3584  <= TRANSPORT DIN(4)  ;
and2_3153: n_3585 <=  n_3586  AND n_3587;
delay_3154: n_3586  <= TRANSPORT a_N1198_aOUT  ;
delay_3155: n_3587  <= TRANSPORT a_N2027_aQ  ;
and1_3156: n_3588 <=  gnd;
inv_3157: n_3589  <= TRANSPORT NOT nTXC  ;
filter_3158: FILTER_a8251
    PORT MAP (IN1 => n_3589, Y => a_N2027_aCLK);
dff_3159: DFF_a8251
    PORT MAP ( D => a_N2026_aD, CLK => a_N2026_aCLK, CLRN => a_N2026_aCLRN,
          PRN => vcc, Q => a_N2026_aQ);
delay_3160: a_N2026_aCLRN  <= TRANSPORT nRESET  ;
xor2_3161: a_N2026_aD <=  n_3597  XOR n_3604;
or2_3162: n_3597 <=  n_3598  OR n_3601;
and2_3163: n_3598 <=  n_3599  AND n_3600;
delay_3164: n_3599  <= TRANSPORT a_N1197_aOUT  ;
delay_3165: n_3600  <= TRANSPORT DIN(5)  ;
and2_3166: n_3601 <=  n_3602  AND n_3603;
delay_3167: n_3602  <= TRANSPORT a_N1198_aOUT  ;
delay_3168: n_3603  <= TRANSPORT a_N2026_aQ  ;
and1_3169: n_3604 <=  gnd;
inv_3170: n_3605  <= TRANSPORT NOT nTXC  ;
filter_3171: FILTER_a8251
    PORT MAP (IN1 => n_3605, Y => a_N2026_aCLK);
dff_3172: DFF_a8251
    PORT MAP ( D => a_N2025_aD, CLK => a_N2025_aCLK, CLRN => a_N2025_aCLRN,
          PRN => vcc, Q => a_N2025_aQ);
delay_3173: a_N2025_aCLRN  <= TRANSPORT nRESET  ;
xor2_3174: a_N2025_aD <=  n_3613  XOR n_3622;
or2_3175: n_3613 <=  n_3614  OR n_3618;
and3_3176: n_3614 <=  n_3615  AND n_3616  AND n_3617;
delay_3177: n_3615  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_3178: n_3616  <= TRANSPORT a_N489_aNOT_aOUT  ;
delay_3179: n_3617  <= TRANSPORT DIN(6)  ;
and3_3180: n_3618 <=  n_3619  AND n_3620  AND n_3621;
delay_3181: n_3619  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_3182: n_3620  <= TRANSPORT NOT a_N489_aNOT_aOUT  ;
delay_3183: n_3621  <= TRANSPORT a_N2025_aQ  ;
and1_3184: n_3622 <=  gnd;
inv_3185: n_3623  <= TRANSPORT NOT nTXC  ;
filter_3186: FILTER_a8251
    PORT MAP (IN1 => n_3623, Y => a_N2025_aCLK);
dff_3187: DFF_a8251
    PORT MAP ( D => a_N2024_aD, CLK => a_N2024_aCLK, CLRN => a_N2024_aCLRN,
          PRN => vcc, Q => a_N2024_aQ);
delay_3188: a_N2024_aCLRN  <= TRANSPORT nRESET  ;
xor2_3189: a_N2024_aD <=  n_3631  XOR n_3640;
or2_3190: n_3631 <=  n_3632  OR n_3636;
and3_3191: n_3632 <=  n_3633  AND n_3634  AND n_3635;
delay_3192: n_3633  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_3193: n_3634  <= TRANSPORT a_N489_aNOT_aOUT  ;
delay_3194: n_3635  <= TRANSPORT DIN(7)  ;
and3_3195: n_3636 <=  n_3637  AND n_3638  AND n_3639;
delay_3196: n_3637  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_3197: n_3638  <= TRANSPORT NOT a_N489_aNOT_aOUT  ;
delay_3198: n_3639  <= TRANSPORT a_N2024_aQ  ;
and1_3199: n_3640 <=  gnd;
inv_3200: n_3641  <= TRANSPORT NOT nTXC  ;
filter_3201: FILTER_a8251
    PORT MAP (IN1 => n_3641, Y => a_N2024_aCLK);
delay_3202: a_N1165_aOUT  <= TRANSPORT a_N1165_aIN  ;
xor2_3203: a_N1165_aIN <=  n_3644  XOR n_3648;
or1_3204: n_3644 <=  n_3645;
and2_3205: n_3645 <=  n_3646  AND n_3647;
delay_3206: n_3646  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3207: n_3647  <= TRANSPORT nRESET  ;
and1_3208: n_3648 <=  gnd;
delay_3209: a_N608_aOUT  <= TRANSPORT a_N608_aIN  ;
xor2_3210: a_N608_aIN <=  n_3651  XOR n_3655;
or1_3211: n_3651 <=  n_3652;
and2_3212: n_3652 <=  n_3653  AND n_3654;
inv_3213: n_3653  <= TRANSPORT NOT a_N1035_aOUT  ;
delay_3214: n_3654  <= TRANSPORT a_N1165_aOUT  ;
and1_3215: n_3655 <=  gnd;
delay_3216: a_LC5_B5_aOUT  <= TRANSPORT a_LC5_B5_aIN  ;
xor2_3217: a_LC5_B5_aIN <=  n_3658  XOR n_3663;
or1_3218: n_3658 <=  n_3659;
and3_3219: n_3659 <=  n_3660  AND n_3661  AND n_3662;
delay_3220: n_3660  <= TRANSPORT a_N1165_aOUT  ;
inv_3221: n_3661  <= TRANSPORT NOT a_N1757_aQ  ;
delay_3222: n_3662  <= TRANSPORT a_N1756_aQ  ;
and1_3223: n_3663 <=  gnd;
delay_3224: a_N120_aOUT  <= TRANSPORT a_N120_aIN  ;
xor2_3225: a_N120_aIN <=  n_3666  XOR n_3670;
or1_3226: n_3666 <=  n_3667;
and2_3227: n_3667 <=  n_3668  AND n_3669;
delay_3228: n_3668  <= TRANSPORT a_N1189_aOUT  ;
delay_3229: n_3669  <= TRANSPORT DIN(1)  ;
and1_3230: n_3670 <=  gnd;
dff_3231: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F1_G_aD, CLK => a_SSYNC1_F1_G_aCLK, CLRN => a_SSYNC1_F1_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F1_G_aQ);
delay_3232: a_SSYNC1_F1_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3233: a_SSYNC1_F1_G_aD <=  n_3678  XOR n_3685;
or2_3234: n_3678 <=  n_3679  OR n_3682;
and2_3235: n_3679 <=  n_3680  AND n_3681;
delay_3236: n_3680  <= TRANSPORT a_N608_aOUT  ;
delay_3237: n_3681  <= TRANSPORT a_SSYNC1_F1_G_aQ  ;
and2_3238: n_3682 <=  n_3683  AND n_3684;
delay_3239: n_3683  <= TRANSPORT a_LC5_B5_aOUT  ;
delay_3240: n_3684  <= TRANSPORT a_N120_aOUT  ;
and1_3241: n_3685 <=  gnd;
delay_3242: n_3686  <= TRANSPORT CLK  ;
filter_3243: FILTER_a8251
    PORT MAP (IN1 => n_3686, Y => a_SSYNC1_F1_G_aCLK);
delay_3244: a_N1168_aNOT_aOUT  <= TRANSPORT a_N1168_aNOT_aIN  ;
xor2_3245: a_N1168_aNOT_aIN <=  n_3690  XOR n_3695;
or2_3246: n_3690 <=  n_3691  OR n_3693;
and1_3247: n_3691 <=  n_3692;
inv_3248: n_3692  <= TRANSPORT NOT a_N1756_aQ  ;
and1_3249: n_3693 <=  n_3694;
inv_3250: n_3694  <= TRANSPORT NOT a_N1757_aQ  ;
and1_3251: n_3695 <=  gnd;
delay_3252: a_N1116_aNOT_aOUT  <= TRANSPORT a_N1116_aNOT_aIN  ;
xor2_3253: a_N1116_aNOT_aIN <=  n_3698  XOR n_3703;
or2_3254: n_3698 <=  n_3699  OR n_3701;
and1_3255: n_3699 <=  n_3700;
delay_3256: n_3700  <= TRANSPORT a_N1168_aNOT_aOUT  ;
and1_3257: n_3701 <=  n_3702;
inv_3258: n_3702  <= TRANSPORT NOT a_N124_aOUT  ;
and1_3259: n_3703 <=  gnd;
delay_3260: a_N718_aOUT  <= TRANSPORT a_N718_aIN  ;
xor2_3261: a_N718_aIN <=  n_3706  XOR n_3711;
or1_3262: n_3706 <=  n_3707;
and3_3263: n_3707 <=  n_3708  AND n_3709  AND n_3710;
delay_3264: n_3708  <= TRANSPORT a_N1189_aOUT  ;
inv_3265: n_3709  <= TRANSPORT NOT a_N1168_aNOT_aOUT  ;
delay_3266: n_3710  <= TRANSPORT DIN(1)  ;
and1_3267: n_3711 <=  gnd;
dff_3268: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F1_G_aD, CLK => a_SSYNC2_F1_G_aCLK, CLRN => a_SSYNC2_F1_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F1_G_aQ);
delay_3269: a_SSYNC2_F1_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3270: a_SSYNC2_F1_G_aD <=  n_3719  XOR n_3727;
or2_3271: n_3719 <=  n_3720  OR n_3724;
and3_3272: n_3720 <=  n_3721  AND n_3722  AND n_3723;
delay_3273: n_3721  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3274: n_3722  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3275: n_3723  <= TRANSPORT a_SSYNC2_F1_G_aQ  ;
and2_3276: n_3724 <=  n_3725  AND n_3726;
delay_3277: n_3725  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3278: n_3726  <= TRANSPORT a_N718_aOUT  ;
and1_3279: n_3727 <=  gnd;
delay_3280: n_3728  <= TRANSPORT CLK  ;
filter_3281: FILTER_a8251
    PORT MAP (IN1 => n_3728, Y => a_SSYNC2_F1_G_aCLK);
delay_3282: a_N723_aOUT  <= TRANSPORT a_N723_aIN  ;
xor2_3283: a_N723_aIN <=  n_3732  XOR n_3738;
or1_3284: n_3732 <=  n_3733;
and4_3285: n_3733 <=  n_3734  AND n_3735  AND n_3736  AND n_3737;
delay_3286: n_3734  <= TRANSPORT a_N1189_aOUT  ;
delay_3287: n_3735  <= TRANSPORT DIN(2)  ;
delay_3288: n_3736  <= TRANSPORT a_N1757_aQ  ;
delay_3289: n_3737  <= TRANSPORT a_N1756_aQ  ;
and1_3290: n_3738 <=  gnd;
dff_3291: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F2_G_aD, CLK => a_SSYNC2_F2_G_aCLK, CLRN => a_SSYNC2_F2_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F2_G_aQ);
delay_3292: a_SSYNC2_F2_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3293: a_SSYNC2_F2_G_aD <=  n_3745  XOR n_3753;
or2_3294: n_3745 <=  n_3746  OR n_3750;
and3_3295: n_3746 <=  n_3747  AND n_3748  AND n_3749;
delay_3296: n_3747  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3297: n_3748  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3298: n_3749  <= TRANSPORT a_SSYNC2_F2_G_aQ  ;
and2_3299: n_3750 <=  n_3751  AND n_3752;
delay_3300: n_3751  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3301: n_3752  <= TRANSPORT a_N723_aOUT  ;
and1_3302: n_3753 <=  gnd;
delay_3303: n_3754  <= TRANSPORT CLK  ;
filter_3304: FILTER_a8251
    PORT MAP (IN1 => n_3754, Y => a_SSYNC2_F2_G_aCLK);
delay_3305: a_N103_aOUT  <= TRANSPORT a_N103_aIN  ;
xor2_3306: a_N103_aIN <=  n_3758  XOR n_3763;
or1_3307: n_3758 <=  n_3759;
and3_3308: n_3759 <=  n_3760  AND n_3761  AND n_3762;
delay_3309: n_3760  <= TRANSPORT a_N1189_aOUT  ;
delay_3310: n_3761  <= TRANSPORT DIN(2)  ;
delay_3311: n_3762  <= TRANSPORT a_N1756_aQ  ;
and1_3312: n_3763 <=  gnd;
dff_3313: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F2_G_aD, CLK => a_SSYNC1_F2_G_aCLK, CLRN => a_SSYNC1_F2_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F2_G_aQ);
delay_3314: a_SSYNC1_F2_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3315: a_SSYNC1_F2_G_aD <=  n_3770  XOR n_3777;
or2_3316: n_3770 <=  n_3771  OR n_3774;
and2_3317: n_3771 <=  n_3772  AND n_3773;
delay_3318: n_3772  <= TRANSPORT a_N608_aOUT  ;
delay_3319: n_3773  <= TRANSPORT a_SSYNC1_F2_G_aQ  ;
and2_3320: n_3774 <=  n_3775  AND n_3776;
delay_3321: n_3775  <= TRANSPORT a_LC5_B5_aOUT  ;
delay_3322: n_3776  <= TRANSPORT a_N103_aOUT  ;
and1_3323: n_3777 <=  gnd;
delay_3324: n_3778  <= TRANSPORT CLK  ;
filter_3325: FILTER_a8251
    PORT MAP (IN1 => n_3778, Y => a_SSYNC1_F2_G_aCLK);
delay_3326: a_LC4_C5_aOUT  <= TRANSPORT a_LC4_C5_aIN  ;
xor2_3327: a_LC4_C5_aIN <=  n_3782  XOR n_3787;
or1_3328: n_3782 <=  n_3783;
and3_3329: n_3783 <=  n_3784  AND n_3785  AND n_3786;
delay_3330: n_3784  <= TRANSPORT a_N1189_aOUT  ;
inv_3331: n_3785  <= TRANSPORT NOT a_N1168_aNOT_aOUT  ;
delay_3332: n_3786  <= TRANSPORT DIN(3)  ;
and1_3333: n_3787 <=  gnd;
dff_3334: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F3_G_aD, CLK => a_SSYNC2_F3_G_aCLK, CLRN => a_SSYNC2_F3_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F3_G_aQ);
delay_3335: a_SSYNC2_F3_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3336: a_SSYNC2_F3_G_aD <=  n_3794  XOR n_3802;
or2_3337: n_3794 <=  n_3795  OR n_3799;
and3_3338: n_3795 <=  n_3796  AND n_3797  AND n_3798;
delay_3339: n_3796  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3340: n_3797  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3341: n_3798  <= TRANSPORT a_SSYNC2_F3_G_aQ  ;
and2_3342: n_3799 <=  n_3800  AND n_3801;
delay_3343: n_3800  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3344: n_3801  <= TRANSPORT a_LC4_C5_aOUT  ;
and1_3345: n_3802 <=  gnd;
delay_3346: n_3803  <= TRANSPORT CLK  ;
filter_3347: FILTER_a8251
    PORT MAP (IN1 => n_3803, Y => a_SSYNC2_F3_G_aCLK);
delay_3348: a_N607_aOUT  <= TRANSPORT a_N607_aIN  ;
xor2_3349: a_N607_aIN <=  n_3806  XOR n_3812;
or1_3350: n_3806 <=  n_3807;
and4_3351: n_3807 <=  n_3808  AND n_3809  AND n_3810  AND n_3811;
delay_3352: n_3808  <= TRANSPORT a_N1189_aOUT  ;
delay_3353: n_3809  <= TRANSPORT a_N1165_aOUT  ;
inv_3354: n_3810  <= TRANSPORT NOT a_N1757_aQ  ;
delay_3355: n_3811  <= TRANSPORT DIN(3)  ;
and1_3356: n_3812 <=  gnd;
dff_3357: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F3_G_aD, CLK => a_SSYNC1_F3_G_aCLK, CLRN => a_SSYNC1_F3_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F3_G_aQ);
delay_3358: a_SSYNC1_F3_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3359: a_SSYNC1_F3_G_aD <=  n_3819  XOR n_3826;
or2_3360: n_3819 <=  n_3820  OR n_3823;
and2_3361: n_3820 <=  n_3821  AND n_3822;
delay_3362: n_3821  <= TRANSPORT a_N608_aOUT  ;
delay_3363: n_3822  <= TRANSPORT a_SSYNC1_F3_G_aQ  ;
and2_3364: n_3823 <=  n_3824  AND n_3825;
delay_3365: n_3824  <= TRANSPORT a_N607_aOUT  ;
delay_3366: n_3825  <= TRANSPORT a_N1756_aQ  ;
and1_3367: n_3826 <=  gnd;
delay_3368: n_3827  <= TRANSPORT CLK  ;
filter_3369: FILTER_a8251
    PORT MAP (IN1 => n_3827, Y => a_SSYNC1_F3_G_aCLK);
dff_3370: DFF_a8251
    PORT MAP ( D => a_N363_aD, CLK => a_N363_aCLK, CLRN => a_N363_aCLRN, PRN => vcc,
          Q => a_N363_aQ);
delay_3371: a_N363_aCLRN  <= TRANSPORT nRESET  ;
xor2_3372: a_N363_aD <=  n_3835  XOR n_3847;
or3_3373: n_3835 <=  n_3836  OR n_3840  OR n_3844;
and3_3374: n_3836 <=  n_3837  AND n_3838  AND n_3839;
inv_3375: n_3837  <= TRANSPORT NOT a_LC4_B6_aNOT_aOUT  ;
delay_3376: n_3838  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_3377: n_3839  <= TRANSPORT NOT a_N363_aQ  ;
and3_3378: n_3840 <=  n_3841  AND n_3842  AND n_3843;
delay_3379: n_3841  <= TRANSPORT a_LC4_B6_aNOT_aOUT  ;
delay_3380: n_3842  <= TRANSPORT a_LC4_B10_aOUT  ;
delay_3381: n_3843  <= TRANSPORT a_N363_aQ  ;
and2_3382: n_3844 <=  n_3845  AND n_3846;
delay_3383: n_3845  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_3384: n_3846  <= TRANSPORT a_N363_aQ  ;
and1_3385: n_3847 <=  gnd;
inv_3386: n_3848  <= TRANSPORT NOT nTXC  ;
filter_3387: FILTER_a8251
    PORT MAP (IN1 => n_3848, Y => a_N363_aCLK);
dff_3388: DFF_a8251
    PORT MAP ( D => a_N362_aD, CLK => a_N362_aCLK, CLRN => a_N362_aCLRN, PRN => vcc,
          Q => a_N362_aQ);
delay_3389: a_N362_aCLRN  <= TRANSPORT nRESET  ;
xor2_3390: a_N362_aD <=  n_3856  XOR n_3868;
or3_3391: n_3856 <=  n_3857  OR n_3861  OR n_3865;
and3_3392: n_3857 <=  n_3858  AND n_3859  AND n_3860;
delay_3393: n_3858  <= TRANSPORT a_LC7_B6_aNOT_aOUT  ;
delay_3394: n_3859  <= TRANSPORT a_LC4_B10_aOUT  ;
delay_3395: n_3860  <= TRANSPORT a_N362_aQ  ;
and3_3396: n_3861 <=  n_3862  AND n_3863  AND n_3864;
inv_3397: n_3862  <= TRANSPORT NOT a_LC7_B6_aNOT_aOUT  ;
delay_3398: n_3863  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_3399: n_3864  <= TRANSPORT NOT a_N362_aQ  ;
and2_3400: n_3865 <=  n_3866  AND n_3867;
delay_3401: n_3866  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_3402: n_3867  <= TRANSPORT a_N362_aQ  ;
and1_3403: n_3868 <=  gnd;
inv_3404: n_3869  <= TRANSPORT NOT nTXC  ;
filter_3405: FILTER_a8251
    PORT MAP (IN1 => n_3869, Y => a_N362_aCLK);
delay_3406: a_LC8_B1_aOUT  <= TRANSPORT a_LC8_B1_aIN  ;
xor2_3407: a_LC8_B1_aIN <=  n_3873  XOR n_3878;
or1_3408: n_3873 <=  n_3874;
and3_3409: n_3874 <=  n_3875  AND n_3876  AND n_3877;
inv_3410: n_3875  <= TRANSPORT NOT a_LC7_B6_aNOT_aOUT  ;
delay_3411: n_3876  <= TRANSPORT a_N362_aQ  ;
delay_3412: n_3877  <= TRANSPORT a_N361_aQ  ;
and1_3413: n_3878 <=  gnd;
dff_3414: DFF_a8251
    PORT MAP ( D => a_N360_aD, CLK => a_N360_aCLK, CLRN => a_N360_aCLRN, PRN => vcc,
          Q => a_N360_aQ);
delay_3415: a_N360_aCLRN  <= TRANSPORT nRESET  ;
xor2_3416: a_N360_aD <=  n_3885  XOR n_3897;
or3_3417: n_3885 <=  n_3886  OR n_3890  OR n_3894;
and3_3418: n_3886 <=  n_3887  AND n_3888  AND n_3889;
delay_3419: n_3887  <= TRANSPORT a_LC4_B10_aOUT  ;
delay_3420: n_3888  <= TRANSPORT a_LC8_B1_aOUT  ;
inv_3421: n_3889  <= TRANSPORT NOT a_N360_aQ  ;
and3_3422: n_3890 <=  n_3891  AND n_3892  AND n_3893;
delay_3423: n_3891  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_3424: n_3892  <= TRANSPORT NOT a_LC8_B1_aOUT  ;
delay_3425: n_3893  <= TRANSPORT a_N360_aQ  ;
and2_3426: n_3894 <=  n_3895  AND n_3896;
delay_3427: n_3895  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_3428: n_3896  <= TRANSPORT a_N360_aQ  ;
and1_3429: n_3897 <=  gnd;
inv_3430: n_3898  <= TRANSPORT NOT nTXC  ;
filter_3431: FILTER_a8251
    PORT MAP (IN1 => n_3898, Y => a_N360_aCLK);
delay_3432: a_LC7_B1_aOUT  <= TRANSPORT a_LC7_B1_aIN  ;
xor2_3433: a_LC7_B1_aIN <=  n_3902  XOR n_3906;
or1_3434: n_3902 <=  n_3903;
and2_3435: n_3903 <=  n_3904  AND n_3905;
inv_3436: n_3904  <= TRANSPORT NOT a_LC7_B6_aNOT_aOUT  ;
delay_3437: n_3905  <= TRANSPORT a_N362_aQ  ;
and1_3438: n_3906 <=  gnd;
dff_3439: DFF_a8251
    PORT MAP ( D => a_N361_aD, CLK => a_N361_aCLK, CLRN => a_N361_aCLRN, PRN => vcc,
          Q => a_N361_aQ);
delay_3440: a_N361_aCLRN  <= TRANSPORT nRESET  ;
xor2_3441: a_N361_aD <=  n_3913  XOR n_3925;
or3_3442: n_3913 <=  n_3914  OR n_3918  OR n_3922;
and3_3443: n_3914 <=  n_3915  AND n_3916  AND n_3917;
delay_3444: n_3915  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_3445: n_3916  <= TRANSPORT NOT a_LC7_B1_aOUT  ;
delay_3446: n_3917  <= TRANSPORT a_N361_aQ  ;
and3_3447: n_3918 <=  n_3919  AND n_3920  AND n_3921;
delay_3448: n_3919  <= TRANSPORT a_LC4_B10_aOUT  ;
delay_3449: n_3920  <= TRANSPORT a_LC7_B1_aOUT  ;
inv_3450: n_3921  <= TRANSPORT NOT a_N361_aQ  ;
and2_3451: n_3922 <=  n_3923  AND n_3924;
delay_3452: n_3923  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_3453: n_3924  <= TRANSPORT a_N361_aQ  ;
and1_3454: n_3925 <=  gnd;
inv_3455: n_3926  <= TRANSPORT NOT nTXC  ;
filter_3456: FILTER_a8251
    PORT MAP (IN1 => n_3926, Y => a_N361_aCLK);
delay_3457: a_N234_aNOT_aOUT  <= TRANSPORT a_N234_aNOT_aIN  ;
xor2_3458: a_N234_aNOT_aIN <=  n_3930  XOR n_3936;
or1_3459: n_3930 <=  n_3931;
and4_3460: n_3931 <=  n_3932  AND n_3933  AND n_3934  AND n_3935;
delay_3461: n_3932  <= TRANSPORT a_N124_aOUT  ;
delay_3462: n_3933  <= TRANSPORT a_N1165_aOUT  ;
inv_3463: n_3934  <= TRANSPORT NOT a_N1168_aNOT_aOUT  ;
delay_3464: n_3935  <= TRANSPORT DIN(6)  ;
and1_3465: n_3936 <=  gnd;
dff_3466: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F6_G_aD, CLK => a_SSYNC2_F6_G_aCLK, CLRN => a_SSYNC2_F6_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F6_G_aQ);
delay_3467: a_SSYNC2_F6_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3468: a_SSYNC2_F6_G_aD <=  n_3943  XOR n_3950;
or2_3469: n_3943 <=  n_3944  OR n_3946;
and1_3470: n_3944 <=  n_3945;
delay_3471: n_3945  <= TRANSPORT a_N234_aNOT_aOUT  ;
and3_3472: n_3946 <=  n_3947  AND n_3948  AND n_3949;
delay_3473: n_3947  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3474: n_3948  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3475: n_3949  <= TRANSPORT a_SSYNC2_F6_G_aQ  ;
and1_3476: n_3950 <=  gnd;
delay_3477: n_3951  <= TRANSPORT CLK  ;
filter_3478: FILTER_a8251
    PORT MAP (IN1 => n_3951, Y => a_SSYNC2_F6_G_aCLK);
dff_3479: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F7_G_aD, CLK => a_SSYNC2_F7_G_aCLK, CLRN => a_SSYNC2_F7_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F7_G_aQ);
delay_3480: a_SSYNC2_F7_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3481: a_SSYNC2_F7_G_aD <=  n_3959  XOR n_3968;
or2_3482: n_3959 <=  n_3960  OR n_3964;
and3_3483: n_3960 <=  n_3961  AND n_3962  AND n_3963;
delay_3484: n_3961  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3485: n_3962  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3486: n_3963  <= TRANSPORT a_SSYNC2_F7_G_aQ  ;
and3_3487: n_3964 <=  n_3965  AND n_3966  AND n_3967;
delay_3488: n_3965  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_3489: n_3966  <= TRANSPORT NOT a_N1116_aNOT_aOUT  ;
delay_3490: n_3967  <= TRANSPORT DIN(7)  ;
and1_3491: n_3968 <=  gnd;
delay_3492: n_3969  <= TRANSPORT CLK  ;
filter_3493: FILTER_a8251
    PORT MAP (IN1 => n_3969, Y => a_SSYNC2_F7_G_aCLK);
delay_3494: a_N233_aNOT_aOUT  <= TRANSPORT a_N233_aNOT_aIN  ;
xor2_3495: a_N233_aNOT_aIN <=  n_3973  XOR n_3979;
or1_3496: n_3973 <=  n_3974;
and4_3497: n_3974 <=  n_3975  AND n_3976  AND n_3977  AND n_3978;
delay_3498: n_3975  <= TRANSPORT a_N124_aOUT  ;
delay_3499: n_3976  <= TRANSPORT a_N1165_aOUT  ;
inv_3500: n_3977  <= TRANSPORT NOT a_N1168_aNOT_aOUT  ;
delay_3501: n_3978  <= TRANSPORT DIN(5)  ;
and1_3502: n_3979 <=  gnd;
dff_3503: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F5_G_aD, CLK => a_SSYNC2_F5_G_aCLK, CLRN => a_SSYNC2_F5_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F5_G_aQ);
delay_3504: a_SSYNC2_F5_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3505: a_SSYNC2_F5_G_aD <=  n_3986  XOR n_3993;
or2_3506: n_3986 <=  n_3987  OR n_3989;
and1_3507: n_3987 <=  n_3988;
delay_3508: n_3988  <= TRANSPORT a_N233_aNOT_aOUT  ;
and3_3509: n_3989 <=  n_3990  AND n_3991  AND n_3992;
delay_3510: n_3990  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3511: n_3991  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3512: n_3992  <= TRANSPORT a_SSYNC2_F5_G_aQ  ;
and1_3513: n_3993 <=  gnd;
delay_3514: n_3994  <= TRANSPORT CLK  ;
filter_3515: FILTER_a8251
    PORT MAP (IN1 => n_3994, Y => a_SSYNC2_F5_G_aCLK);
dff_3516: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F4_G_aD, CLK => a_SSYNC2_F4_G_aCLK, CLRN => a_SSYNC2_F4_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F4_G_aQ);
delay_3517: a_SSYNC2_F4_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_3518: a_SSYNC2_F4_G_aD <=  n_4002  XOR n_4011;
or2_3519: n_4002 <=  n_4003  OR n_4007;
and3_3520: n_4003 <=  n_4004  AND n_4005  AND n_4006;
delay_3521: n_4004  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_3522: n_4005  <= TRANSPORT NOT a_N1116_aNOT_aOUT  ;
delay_3523: n_4006  <= TRANSPORT DIN(4)  ;
and3_3524: n_4007 <=  n_4008  AND n_4009  AND n_4010;
delay_3525: n_4008  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_3526: n_4009  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_3527: n_4010  <= TRANSPORT a_SSYNC2_F4_G_aQ  ;
and1_3528: n_4011 <=  gnd;
delay_3529: n_4012  <= TRANSPORT CLK  ;
filter_3530: FILTER_a8251
    PORT MAP (IN1 => n_4012, Y => a_SSYNC2_F4_G_aCLK);
delay_3531: a_N1120_aNOT_aOUT  <= TRANSPORT a_N1120_aNOT_aIN  ;
xor2_3532: a_N1120_aNOT_aIN <=  n_4015  XOR n_4022;
or2_3533: n_4015 <=  n_4016  OR n_4019;
and1_3534: n_4016 <=  n_4017;
delay_3535: n_4017  <= TRANSPORT a_N1902_aQ  ;
and1_3536: n_4019 <=  n_4020;
inv_3537: n_4020  <= TRANSPORT NOT a_N1901_aQ  ;
and1_3538: n_4022 <=  gnd;
delay_3539: a_N1052_aOUT  <= TRANSPORT a_N1052_aIN  ;
xor2_3540: a_N1052_aIN <=  n_4025  XOR n_4029;
or1_3541: n_4025 <=  n_4026;
and2_3542: n_4026 <=  n_4027  AND n_4028;
delay_3543: n_4027  <= TRANSPORT a_N1138_aOUT  ;
delay_3544: n_4028  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3545: n_4029 <=  gnd;
delay_3546: a_N1177_aOUT  <= TRANSPORT a_N1177_aIN  ;
xor2_3547: a_N1177_aIN <=  n_4032  XOR n_4043;
or2_3548: n_4032 <=  n_4033  OR n_4039;
and3_3549: n_4033 <=  n_4034  AND n_4036  AND n_4038;
inv_3550: n_4034  <= TRANSPORT NOT a_N1555_aQ  ;
delay_3551: n_4036  <= TRANSPORT a_N1556_aQ  ;
inv_3552: n_4038  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and3_3553: n_4039 <=  n_4040  AND n_4041  AND n_4042;
delay_3554: n_4040  <= TRANSPORT a_N1555_aQ  ;
inv_3555: n_4041  <= TRANSPORT NOT a_N1556_aQ  ;
inv_3556: n_4042  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_3557: n_4043 <=  gnd;
delay_3558: a_N420_aOUT  <= TRANSPORT a_N420_aIN  ;
xor2_3559: a_N420_aIN <=  n_4046  XOR n_4055;
or4_3560: n_4046 <=  n_4047  OR n_4049  OR n_4051  OR n_4053;
and1_3561: n_4047 <=  n_4048;
inv_3562: n_4048  <= TRANSPORT NOT a_N1052_aOUT  ;
and1_3563: n_4049 <=  n_4050;
inv_3564: n_4050  <= TRANSPORT NOT a_N1177_aOUT  ;
and1_3565: n_4051 <=  n_4052;
inv_3566: n_4052  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_3567: n_4053 <=  n_4054;
delay_3568: n_4054  <= TRANSPORT a_N83_aOUT  ;
and1_3569: n_4055 <=  gnd;
delay_3570: a_LC3_A1_aOUT  <= TRANSPORT a_LC3_A1_aIN  ;
xor2_3571: a_LC3_A1_aIN <=  n_4058  XOR n_4069;
or2_3572: n_4058 <=  n_4059  OR n_4064;
and4_3573: n_4059 <=  n_4060  AND n_4061  AND n_4062  AND n_4063;
inv_3574: n_4060  <= TRANSPORT NOT a_N83_aOUT  ;
inv_3575: n_4061  <= TRANSPORT NOT a_N1555_aQ  ;
delay_3576: n_4062  <= TRANSPORT a_N1556_aQ  ;
inv_3577: n_4063  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and4_3578: n_4064 <=  n_4065  AND n_4066  AND n_4067  AND n_4068;
inv_3579: n_4065  <= TRANSPORT NOT a_N83_aOUT  ;
delay_3580: n_4066  <= TRANSPORT a_N1555_aQ  ;
inv_3581: n_4067  <= TRANSPORT NOT a_N1556_aQ  ;
inv_3582: n_4068  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_3583: n_4069 <=  gnd;
delay_3584: a_LC4_A1_aOUT  <= TRANSPORT a_LC4_A1_aIN  ;
xor2_3585: a_LC4_A1_aIN <=  n_4072  XOR n_4083;
or2_3586: n_4072 <=  n_4073  OR n_4078;
and4_3587: n_4073 <=  n_4074  AND n_4075  AND n_4076  AND n_4077;
delay_3588: n_4074  <= TRANSPORT a_LC3_A1_aOUT  ;
delay_3589: n_4075  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
delay_3590: n_4076  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
inv_3591: n_4077  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and4_3592: n_4078 <=  n_4079  AND n_4080  AND n_4081  AND n_4082;
delay_3593: n_4079  <= TRANSPORT a_LC3_A1_aOUT  ;
delay_3594: n_4080  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_3595: n_4081  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
delay_3596: n_4082  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3597: n_4083 <=  gnd;
delay_3598: a_N1050_aOUT  <= TRANSPORT a_N1050_aIN  ;
xor2_3599: a_N1050_aIN <=  n_4086  XOR n_4091;
or1_3600: n_4086 <=  n_4087;
and3_3601: n_4087 <=  n_4088  AND n_4089  AND n_4090;
inv_3602: n_4088  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
delay_3603: n_4089  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
delay_3604: n_4090  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3605: n_4091 <=  gnd;
delay_3606: a_N1187_aOUT  <= TRANSPORT a_N1187_aIN  ;
xor2_3607: a_N1187_aIN <=  n_4094  XOR n_4098;
or1_3608: n_4094 <=  n_4095;
and2_3609: n_4095 <=  n_4096  AND n_4097;
inv_3610: n_4096  <= TRANSPORT NOT a_N83_aOUT  ;
inv_3611: n_4097  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_3612: n_4098 <=  gnd;
delay_3613: a_LC1_A15_aOUT  <= TRANSPORT a_LC1_A15_aIN  ;
xor2_3614: a_LC1_A15_aIN <=  n_4101  XOR n_4112;
or4_3615: n_4101 <=  n_4102  OR n_4104  OR n_4107  OR n_4110;
and1_3616: n_4102 <=  n_4103;
delay_3617: n_4103  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and2_3618: n_4104 <=  n_4105  AND n_4106;
delay_3619: n_4105  <= TRANSPORT a_N1555_aQ  ;
delay_3620: n_4106  <= TRANSPORT a_N1556_aQ  ;
and2_3621: n_4107 <=  n_4108  AND n_4109;
inv_3622: n_4108  <= TRANSPORT NOT a_N1555_aQ  ;
inv_3623: n_4109  <= TRANSPORT NOT a_N1556_aQ  ;
and1_3624: n_4110 <=  n_4111;
inv_3625: n_4111  <= TRANSPORT NOT a_N1187_aOUT  ;
and1_3626: n_4112 <=  gnd;
delay_3627: a_N676_aOUT  <= TRANSPORT a_N676_aIN  ;
xor2_3628: a_N676_aIN <=  n_4115  XOR n_4124;
or2_3629: n_4115 <=  n_4116  OR n_4120;
and3_3630: n_4116 <=  n_4117  AND n_4118  AND n_4119;
delay_3631: n_4117  <= TRANSPORT a_N1187_aOUT  ;
inv_3632: n_4118  <= TRANSPORT NOT a_N1555_aQ  ;
delay_3633: n_4119  <= TRANSPORT a_N1556_aQ  ;
and3_3634: n_4120 <=  n_4121  AND n_4122  AND n_4123;
delay_3635: n_4121  <= TRANSPORT a_N1187_aOUT  ;
delay_3636: n_4122  <= TRANSPORT a_N1555_aQ  ;
inv_3637: n_4123  <= TRANSPORT NOT a_N1556_aQ  ;
and1_3638: n_4124 <=  gnd;
delay_3639: a_N1135_aNOT_aOUT  <= TRANSPORT a_N1135_aNOT_aIN  ;
xor2_3640: a_N1135_aNOT_aIN <=  n_4127  XOR n_4132;
or2_3641: n_4127 <=  n_4128  OR n_4130;
and1_3642: n_4128 <=  n_4129;
delay_3643: n_4129  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3644: n_4130 <=  n_4131;
inv_3645: n_4131  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and1_3646: n_4132 <=  gnd;
delay_3647: a_LC2_A15_aNOT_aOUT  <= TRANSPORT a_LC2_A15_aNOT_aIN  ;
xor2_3648: a_LC2_A15_aNOT_aIN <=  n_4135  XOR n_4148;
or4_3649: n_4135 <=  n_4136  OR n_4139  OR n_4142  OR n_4145;
and2_3650: n_4136 <=  n_4137  AND n_4138;
inv_3651: n_4137  <= TRANSPORT NOT a_N1050_aOUT  ;
delay_3652: n_4138  <= TRANSPORT a_LC1_A15_aOUT  ;
and2_3653: n_4139 <=  n_4140  AND n_4141;
delay_3654: n_4140  <= TRANSPORT a_LC1_A15_aOUT  ;
inv_3655: n_4141  <= TRANSPORT NOT a_N676_aOUT  ;
and2_3656: n_4142 <=  n_4143  AND n_4144;
inv_3657: n_4143  <= TRANSPORT NOT a_N1050_aOUT  ;
delay_3658: n_4144  <= TRANSPORT a_N1135_aNOT_aOUT  ;
and2_3659: n_4145 <=  n_4146  AND n_4147;
inv_3660: n_4146  <= TRANSPORT NOT a_N676_aOUT  ;
delay_3661: n_4147  <= TRANSPORT a_N1135_aNOT_aOUT  ;
and1_3662: n_4148 <=  gnd;
delay_3663: a_N425_aNOT_aOUT  <= TRANSPORT a_N425_aNOT_aIN  ;
xor2_3664: a_N425_aNOT_aIN <=  n_4151  XOR n_4159;
or3_3665: n_4151 <=  n_4152  OR n_4155  OR n_4157;
and2_3666: n_4152 <=  n_4153  AND n_4154;
delay_3667: n_4153  <= TRANSPORT a_N420_aOUT  ;
delay_3668: n_4154  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_3669: n_4155 <=  n_4156;
delay_3670: n_4156  <= TRANSPORT a_LC4_A1_aOUT  ;
and1_3671: n_4157 <=  n_4158;
inv_3672: n_4158  <= TRANSPORT NOT a_LC2_A15_aNOT_aOUT  ;
and1_3673: n_4159 <=  gnd;
delay_3674: a_N1054_aNOT_aOUT  <= TRANSPORT a_N1054_aNOT_aIN  ;
xor2_3675: a_N1054_aNOT_aIN <=  n_4162  XOR n_4169;
or3_3676: n_4162 <=  n_4163  OR n_4165  OR n_4167;
and1_3677: n_4163 <=  n_4164;
delay_3678: n_4164  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3679: n_4165 <=  n_4166;
delay_3680: n_4166  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_3681: n_4167 <=  n_4168;
delay_3682: n_4168  <= TRANSPORT a_LC1_A15_aOUT  ;
and1_3683: n_4169 <=  gnd;
delay_3684: a_N1049_aNOT_aOUT  <= TRANSPORT a_N1049_aNOT_aIN  ;
xor2_3685: a_N1049_aNOT_aIN <=  n_4172  XOR n_4179;
or3_3686: n_4172 <=  n_4173  OR n_4175  OR n_4177;
and1_3687: n_4173 <=  n_4174;
delay_3688: n_4174  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3689: n_4175 <=  n_4176;
inv_3690: n_4176  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and1_3691: n_4177 <=  n_4178;
delay_3692: n_4178  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and1_3693: n_4179 <=  gnd;
delay_3694: a_LC2_A1_aNOT_aOUT  <= TRANSPORT a_LC2_A1_aNOT_aIN  ;
xor2_3695: a_LC2_A1_aNOT_aIN <=  n_4182  XOR n_4187;
or1_3696: n_4182 <=  n_4183;
and3_3697: n_4183 <=  n_4184  AND n_4185  AND n_4186;
inv_3698: n_4184  <= TRANSPORT NOT a_N83_aOUT  ;
delay_3699: n_4185  <= TRANSPORT a_N1177_aOUT  ;
delay_3700: n_4186  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3701: n_4187 <=  gnd;
delay_3702: a_LC5_A1_aOUT  <= TRANSPORT a_LC5_A1_aIN  ;
xor2_3703: a_LC5_A1_aIN <=  n_4190  XOR n_4197;
or2_3704: n_4190 <=  n_4191  OR n_4194;
and2_3705: n_4191 <=  n_4192  AND n_4193;
delay_3706: n_4192  <= TRANSPORT a_LC3_A1_aOUT  ;
inv_3707: n_4193  <= TRANSPORT NOT a_N1049_aNOT_aOUT  ;
and2_3708: n_4194 <=  n_4195  AND n_4196;
inv_3709: n_4195  <= TRANSPORT NOT a_N1134_aNOT_aOUT  ;
delay_3710: n_4196  <= TRANSPORT a_LC2_A1_aNOT_aOUT  ;
and1_3711: n_4197 <=  gnd;
delay_3712: a_N427_aOUT  <= TRANSPORT a_N427_aIN  ;
xor2_3713: a_N427_aIN <=  n_4200  XOR n_4216;
or4_3714: n_4200 <=  n_4201  OR n_4205  OR n_4208  OR n_4211;
and2_3715: n_4201 <=  n_4202  AND n_4203;
inv_3716: n_4202  <= TRANSPORT NOT a_N425_aNOT_aOUT  ;
delay_3717: n_4203  <= TRANSPORT a_N1170_aQ  ;
and2_3718: n_4205 <=  n_4206  AND n_4207;
inv_3719: n_4206  <= TRANSPORT NOT a_N1054_aNOT_aOUT  ;
delay_3720: n_4207  <= TRANSPORT a_N1170_aQ  ;
and2_3721: n_4208 <=  n_4209  AND n_4210;
delay_3722: n_4209  <= TRANSPORT a_LC5_A1_aOUT  ;
delay_3723: n_4210  <= TRANSPORT a_N1170_aQ  ;
and4_3724: n_4211 <=  n_4212  AND n_4213  AND n_4214  AND n_4215;
delay_3725: n_4212  <= TRANSPORT a_N425_aNOT_aOUT  ;
delay_3726: n_4213  <= TRANSPORT a_N1054_aNOT_aOUT  ;
inv_3727: n_4214  <= TRANSPORT NOT a_LC5_A1_aOUT  ;
inv_3728: n_4215  <= TRANSPORT NOT a_N1170_aQ  ;
and1_3729: n_4216 <=  gnd;
delay_3730: a_N423_aNOT_aOUT  <= TRANSPORT a_N423_aNOT_aIN  ;
xor2_3731: a_N423_aNOT_aIN <=  n_4219  XOR n_4225;
or2_3732: n_4219 <=  n_4220  OR n_4222;
and1_3733: n_4220 <=  n_4221;
delay_3734: n_4221  <= TRANSPORT a_LC4_A1_aOUT  ;
and2_3735: n_4222 <=  n_4223  AND n_4224;
delay_3736: n_4223  <= TRANSPORT a_N420_aOUT  ;
delay_3737: n_4224  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_3738: n_4225 <=  gnd;
delay_3739: a_N428_aOUT  <= TRANSPORT a_N428_aIN  ;
xor2_3740: a_N428_aIN <=  n_4228  XOR n_4236;
or2_3741: n_4228 <=  n_4229  OR n_4232;
and2_3742: n_4229 <=  n_4230  AND n_4231;
delay_3743: n_4230  <= TRANSPORT a_N1054_aNOT_aOUT  ;
delay_3744: n_4231  <= TRANSPORT a_LC5_A1_aOUT  ;
and3_3745: n_4232 <=  n_4233  AND n_4234  AND n_4235;
delay_3746: n_4233  <= TRANSPORT a_LC2_A15_aNOT_aOUT  ;
delay_3747: n_4234  <= TRANSPORT a_N1054_aNOT_aOUT  ;
delay_3748: n_4235  <= TRANSPORT a_N423_aNOT_aOUT  ;
and1_3749: n_4236 <=  gnd;
delay_3750: a_LC2_A12_aOUT  <= TRANSPORT a_LC2_A12_aIN  ;
xor2_3751: a_LC2_A12_aIN <=  n_4239  XOR n_4254;
or4_3752: n_4239 <=  n_4240  OR n_4244  OR n_4248  OR n_4251;
and2_3753: n_4240 <=  n_4241  AND n_4242;
inv_3754: n_4241  <= TRANSPORT NOT a_N420_aOUT  ;
delay_3755: n_4242  <= TRANSPORT a_N1169_aQ  ;
and2_3756: n_4244 <=  n_4245  AND n_4246;
inv_3757: n_4245  <= TRANSPORT NOT a_N420_aOUT  ;
inv_3758: n_4246  <= TRANSPORT NOT a_N1167_aQ  ;
and2_3759: n_4248 <=  n_4249  AND n_4250;
delay_3760: n_4249  <= TRANSPORT a_N420_aOUT  ;
inv_3761: n_4250  <= TRANSPORT NOT a_N1169_aQ  ;
and2_3762: n_4251 <=  n_4252  AND n_4253;
delay_3763: n_4252  <= TRANSPORT a_N420_aOUT  ;
delay_3764: n_4253  <= TRANSPORT a_N1167_aQ  ;
and1_3765: n_4254 <=  gnd;
delay_3766: a_N132_aOUT  <= TRANSPORT a_N132_aIN  ;
xor2_3767: a_N132_aIN <=  n_4257  XOR n_4269;
or4_3768: n_4257 <=  n_4258  OR n_4260  OR n_4264  OR n_4267;
and1_3769: n_4258 <=  n_4259;
delay_3770: n_4259  <= TRANSPORT a_N427_aOUT  ;
and2_3771: n_4260 <=  n_4261  AND n_4262;
inv_3772: n_4261  <= TRANSPORT NOT a_N428_aOUT  ;
delay_3773: n_4262  <= TRANSPORT a_N1171_aQ  ;
and2_3774: n_4264 <=  n_4265  AND n_4266;
delay_3775: n_4265  <= TRANSPORT a_N428_aOUT  ;
inv_3776: n_4266  <= TRANSPORT NOT a_N1171_aQ  ;
and1_3777: n_4267 <=  n_4268;
delay_3778: n_4268  <= TRANSPORT a_LC2_A12_aOUT  ;
and1_3779: n_4269 <=  gnd;
delay_3780: a_N1146_aOUT  <= TRANSPORT a_N1146_aIN  ;
xor2_3781: a_N1146_aIN <=  n_4272  XOR n_4276;
or1_3782: n_4272 <=  n_4273;
and2_3783: n_4273 <=  n_4274  AND n_4275;
inv_3784: n_4274  <= TRANSPORT NOT a_N62_aQ  ;
delay_3785: n_4275  <= TRANSPORT a_N63_aQ  ;
and1_3786: n_4276 <=  gnd;
delay_3787: a_LC1_D2_aNOT_aOUT  <= TRANSPORT a_LC1_D2_aNOT_aIN  ;
xor2_3788: a_LC1_D2_aNOT_aIN <=  n_4279  XOR n_4286;
or3_3789: n_4279 <=  n_4280  OR n_4282  OR n_4284;
and1_3790: n_4280 <=  n_4281;
delay_3791: n_4281  <= TRANSPORT a_N61_aQ  ;
and1_3792: n_4282 <=  n_4283;
inv_3793: n_4283  <= TRANSPORT NOT a_N64_aQ  ;
and1_3794: n_4284 <=  n_4285;
inv_3795: n_4285  <= TRANSPORT NOT a_N1146_aOUT  ;
and1_3796: n_4286 <=  gnd;
delay_3797: a_N1070_aOUT  <= TRANSPORT a_N1070_aIN  ;
xor2_3798: a_N1070_aIN <=  n_4289  XOR n_4295;
or2_3799: n_4289 <=  n_4290  OR n_4293;
and2_3800: n_4290 <=  n_4291  AND n_4292;
delay_3801: n_4291  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_3802: n_4292  <= TRANSPORT a_N132_aOUT  ;
and1_3803: n_4293 <=  n_4294;
delay_3804: n_4294  <= TRANSPORT a_LC1_D2_aNOT_aOUT  ;
and1_3805: n_4295 <=  gnd;
delay_3806: a_LC5_C13_aOUT  <= TRANSPORT a_LC5_C13_aIN  ;
xor2_3807: a_LC5_C13_aIN <=  n_4297  XOR n_4306;
or4_3808: n_4297 <=  n_4298  OR n_4300  OR n_4302  OR n_4304;
and1_3809: n_4298 <=  n_4299;
delay_3810: n_4299  <= TRANSPORT a_N1756_aQ  ;
and1_3811: n_4300 <=  n_4301;
delay_3812: n_4301  <= TRANSPORT a_N1757_aQ  ;
and1_3813: n_4302 <=  n_4303;
inv_3814: n_4303  <= TRANSPORT NOT a_N1754_aQ  ;
and1_3815: n_4304 <=  n_4305;
inv_3816: n_4305  <= TRANSPORT NOT a_N82_aNOT_aOUT  ;
and1_3817: n_4306 <=  gnd;
delay_3818: a_N127_aOUT  <= TRANSPORT a_N127_aIN  ;
xor2_3819: a_N127_aIN <=  n_4309  XOR n_4313;
or1_3820: n_4309 <=  n_4310;
and2_3821: n_4310 <=  n_4311  AND n_4312;
inv_3822: n_4311  <= TRANSPORT NOT a_N64_aQ  ;
inv_3823: n_4312  <= TRANSPORT NOT a_N61_aQ  ;
and1_3824: n_4313 <=  gnd;
delay_3825: a_N1073_aNOT_aOUT  <= TRANSPORT a_N1073_aNOT_aIN  ;
xor2_3826: a_N1073_aNOT_aIN <=  n_4316  XOR n_4325;
or4_3827: n_4316 <=  n_4317  OR n_4319  OR n_4321  OR n_4323;
and1_3828: n_4317 <=  n_4318;
delay_3829: n_4318  <= TRANSPORT a_LC5_C13_aOUT  ;
and1_3830: n_4319 <=  n_4320;
inv_3831: n_4320  <= TRANSPORT NOT a_N127_aOUT  ;
and1_3832: n_4321 <=  n_4322;
delay_3833: n_4322  <= TRANSPORT a_LC2_D19_aOUT  ;
and1_3834: n_4323 <=  n_4324;
delay_3835: n_4324  <= TRANSPORT a_N130_aNOT_aOUT  ;
and1_3836: n_4325 <=  gnd;
delay_3837: a_N1072_aNOT_aOUT  <= TRANSPORT a_N1072_aNOT_aIN  ;
xor2_3838: a_N1072_aNOT_aIN <=  n_4328  XOR n_4337;
or4_3839: n_4328 <=  n_4329  OR n_4331  OR n_4333  OR n_4335;
and1_3840: n_4329 <=  n_4330;
inv_3841: n_4330  <= TRANSPORT NOT a_N63_aQ  ;
and1_3842: n_4331 <=  n_4332;
inv_3843: n_4332  <= TRANSPORT NOT a_N62_aQ  ;
and1_3844: n_4333 <=  n_4334;
delay_3845: n_4334  <= TRANSPORT a_N1152_aNOT_aOUT  ;
and1_3846: n_4335 <=  n_4336;
delay_3847: n_4336  <= TRANSPORT a_N132_aOUT  ;
and1_3848: n_4337 <=  gnd;
delay_3849: a_N1164_aOUT  <= TRANSPORT a_N1164_aIN  ;
xor2_3850: a_N1164_aIN <=  n_4340  XOR n_4344;
or1_3851: n_4340 <=  n_4341;
and2_3852: n_4341 <=  n_4342  AND n_4343;
inv_3853: n_4342  <= TRANSPORT NOT a_N64_aQ  ;
delay_3854: n_4343  <= TRANSPORT a_N61_aQ  ;
and1_3855: n_4344 <=  gnd;
delay_3856: a_N1080_aOUT  <= TRANSPORT a_N1080_aIN  ;
xor2_3857: a_N1080_aIN <=  n_4347  XOR n_4352;
or1_3858: n_4347 <=  n_4348;
and3_3859: n_4348 <=  n_4349  AND n_4350  AND n_4351;
delay_3860: n_4349  <= TRANSPORT a_N1164_aOUT  ;
inv_3861: n_4350  <= TRANSPORT NOT a_N62_aQ  ;
inv_3862: n_4351  <= TRANSPORT NOT a_N63_aQ  ;
and1_3863: n_4352 <=  gnd;
delay_3864: a_LC5_D16_aOUT  <= TRANSPORT a_LC5_D16_aIN  ;
xor2_3865: a_LC5_D16_aIN <=  n_4355  XOR n_4364;
or2_3866: n_4355 <=  n_4356  OR n_4360;
and3_3867: n_4356 <=  n_4357  AND n_4358  AND n_4359;
delay_3868: n_4357  <= TRANSPORT a_N132_aOUT  ;
delay_3869: n_4358  <= TRANSPORT a_N1073_aNOT_aOUT  ;
delay_3870: n_4359  <= TRANSPORT a_N1072_aNOT_aOUT  ;
and3_3871: n_4360 <=  n_4361  AND n_4362  AND n_4363;
delay_3872: n_4361  <= TRANSPORT a_N1073_aNOT_aOUT  ;
delay_3873: n_4362  <= TRANSPORT a_N1072_aNOT_aOUT  ;
inv_3874: n_4363  <= TRANSPORT NOT a_N1080_aOUT  ;
and1_3875: n_4364 <=  gnd;
delay_3876: a_N167_aOUT  <= TRANSPORT a_N167_aIN  ;
xor2_3877: a_N167_aIN <=  n_4367  XOR n_4373;
or1_3878: n_4367 <=  n_4368;
and4_3879: n_4368 <=  n_4369  AND n_4370  AND n_4371  AND n_4372;
delay_3880: n_4369  <= TRANSPORT a_N735_aNOT_aOUT  ;
delay_3881: n_4370  <= TRANSPORT a_N352_aOUT  ;
delay_3882: n_4371  <= TRANSPORT a_N1070_aOUT  ;
delay_3883: n_4372  <= TRANSPORT a_LC5_D16_aOUT  ;
and1_3884: n_4373 <=  gnd;
delay_3885: a_N35_aNOT_aOUT  <= TRANSPORT a_N35_aNOT_aIN  ;
xor2_3886: a_N35_aNOT_aIN <=  n_4376  XOR n_4383;
or2_3887: n_4376 <=  n_4377  OR n_4380;
and2_3888: n_4377 <=  n_4378  AND n_4379;
delay_3889: n_4378  <= TRANSPORT a_N1049_aNOT_aOUT  ;
inv_3890: n_4379  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_3891: n_4380 <=  n_4381  AND n_4382;
delay_3892: n_4381  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_3893: n_4382  <= TRANSPORT a_N1049_aNOT_aOUT  ;
and1_3894: n_4383 <=  gnd;
delay_3895: a_N465_aNOT_aOUT  <= TRANSPORT a_N465_aNOT_aIN  ;
xor2_3896: a_N465_aNOT_aIN <=  n_4386  XOR n_4395;
or2_3897: n_4386 <=  n_4387  OR n_4391;
and2_3898: n_4387 <=  n_4388  AND n_4389;
inv_3899: n_4388  <= TRANSPORT NOT a_N35_aNOT_aOUT  ;
delay_3900: n_4389  <= TRANSPORT a_N1302_aQ  ;
and2_3901: n_4391 <=  n_4392  AND n_4393;
delay_3902: n_4392  <= TRANSPORT a_N35_aNOT_aOUT  ;
delay_3903: n_4393  <= TRANSPORT a_N1301_aQ  ;
and1_3904: n_4395 <=  gnd;
delay_3905: a_N1051_aOUT  <= TRANSPORT a_N1051_aIN  ;
xor2_3906: a_N1051_aIN <=  n_4398  XOR n_4403;
or1_3907: n_4398 <=  n_4399;
and3_3908: n_4399 <=  n_4400  AND n_4401  AND n_4402;
delay_3909: n_4400  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_3910: n_4401  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
inv_3911: n_4402  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_3912: n_4403 <=  gnd;
delay_3913: a_N466_aNOT_aOUT  <= TRANSPORT a_N466_aNOT_aIN  ;
xor2_3914: a_N466_aNOT_aIN <=  n_4406  XOR n_4418;
or3_3915: n_4406 <=  n_4407  OR n_4411  OR n_4415;
and3_3916: n_4407 <=  n_4408  AND n_4409  AND n_4410;
inv_3917: n_4408  <= TRANSPORT NOT a_N1050_aOUT  ;
delay_3918: n_4409  <= TRANSPORT a_N465_aNOT_aOUT  ;
inv_3919: n_4410  <= TRANSPORT NOT a_N1051_aOUT  ;
and2_3920: n_4411 <=  n_4412  AND n_4413;
delay_3921: n_4412  <= TRANSPORT a_N1051_aOUT  ;
delay_3922: n_4413  <= TRANSPORT a_N1303_aQ  ;
and2_3923: n_4415 <=  n_4416  AND n_4417;
delay_3924: n_4416  <= TRANSPORT a_N1050_aOUT  ;
delay_3925: n_4417  <= TRANSPORT a_N1303_aQ  ;
and1_3926: n_4418 <=  gnd;
delay_3927: a_N54_aOUT  <= TRANSPORT a_N54_aIN  ;
xor2_3928: a_N54_aIN <=  n_4421  XOR n_4430;
or2_3929: n_4421 <=  n_4422  OR n_4426;
and3_3930: n_4422 <=  n_4423  AND n_4424  AND n_4425;
delay_3931: n_4423  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
delay_3932: n_4424  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
inv_3933: n_4425  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and3_3934: n_4426 <=  n_4427  AND n_4428  AND n_4429;
delay_3935: n_4427  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_3936: n_4428  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
delay_3937: n_4429  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_3938: n_4430 <=  gnd;
delay_3939: a_N12_aOUT  <= TRANSPORT a_N12_aIN  ;
xor2_3940: a_N12_aIN <=  n_4433  XOR n_4443;
or3_3941: n_4433 <=  n_4434  OR n_4437  OR n_4441;
and2_3942: n_4434 <=  n_4435  AND n_4436;
delay_3943: n_4435  <= TRANSPORT a_N466_aNOT_aOUT  ;
inv_3944: n_4436  <= TRANSPORT NOT a_N54_aOUT  ;
and2_3945: n_4437 <=  n_4438  AND n_4439;
delay_3946: n_4438  <= TRANSPORT a_N54_aOUT  ;
delay_3947: n_4439  <= TRANSPORT a_N1304_aQ  ;
and1_3948: n_4441 <=  n_4442;
delay_3949: n_4442  <= TRANSPORT a_N1052_aOUT  ;
and1_3950: n_4443 <=  gnd;
delay_3951: a_N1102_aNOT_aOUT  <= TRANSPORT a_N1102_aNOT_aIN  ;
xor2_3952: a_N1102_aNOT_aIN <=  n_4445  XOR n_4453;
or2_3953: n_4445 <=  n_4446  OR n_4450;
and2_3954: n_4446 <=  n_4447  AND n_4448;
delay_3955: n_4447  <= TRANSPORT a_N12_aOUT  ;
delay_3956: n_4448  <= TRANSPORT a_N1305_aQ  ;
and2_3957: n_4450 <=  n_4451  AND n_4452;
inv_3958: n_4451  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_3959: n_4452  <= TRANSPORT a_N12_aOUT  ;
and1_3960: n_4453 <=  gnd;
delay_3961: a_N1205_aOUT  <= TRANSPORT a_N1205_aIN  ;
xor2_3962: a_N1205_aIN <=  n_4456  XOR n_4473;
or4_3963: n_4456 <=  n_4457  OR n_4461  OR n_4465  OR n_4469;
and3_3964: n_4457 <=  n_4458  AND n_4459  AND n_4460;
inv_3965: n_4458  <= TRANSPORT NOT a_SSYNC1_F2_G_aQ  ;
delay_3966: n_4459  <= TRANSPORT a_N676_aOUT  ;
delay_3967: n_4460  <= TRANSPORT a_N1102_aNOT_aOUT  ;
and3_3968: n_4461 <=  n_4462  AND n_4463  AND n_4464;
inv_3969: n_4462  <= TRANSPORT NOT a_SSYNC1_F2_G_aQ  ;
inv_3970: n_4463  <= TRANSPORT NOT a_N676_aOUT  ;
delay_3971: n_4464  <= TRANSPORT a_SRXREG_F2_G_aQ  ;
and3_3972: n_4465 <=  n_4466  AND n_4467  AND n_4468;
delay_3973: n_4466  <= TRANSPORT a_SSYNC1_F2_G_aQ  ;
delay_3974: n_4467  <= TRANSPORT a_N676_aOUT  ;
inv_3975: n_4468  <= TRANSPORT NOT a_N1102_aNOT_aOUT  ;
and3_3976: n_4469 <=  n_4470  AND n_4471  AND n_4472;
delay_3977: n_4470  <= TRANSPORT a_SSYNC1_F2_G_aQ  ;
inv_3978: n_4471  <= TRANSPORT NOT a_N676_aOUT  ;
inv_3979: n_4472  <= TRANSPORT NOT a_SRXREG_F2_G_aQ  ;
and1_3980: n_4473 <=  gnd;
delay_3981: a_N1_aOUT  <= TRANSPORT a_N1_aIN  ;
xor2_3982: a_N1_aIN <=  n_4476  XOR n_4485;
or3_3983: n_4476 <=  n_4477  OR n_4480  OR n_4483;
and2_3984: n_4477 <=  n_4478  AND n_4479;
inv_3985: n_4478  <= TRANSPORT NOT a_N35_aNOT_aOUT  ;
delay_3986: n_4479  <= TRANSPORT a_N1303_aQ  ;
and2_3987: n_4480 <=  n_4481  AND n_4482;
delay_3988: n_4481  <= TRANSPORT a_N35_aNOT_aOUT  ;
delay_3989: n_4482  <= TRANSPORT a_N1302_aQ  ;
and1_3990: n_4483 <=  n_4484;
delay_3991: n_4484  <= TRANSPORT a_N1050_aOUT  ;
and1_3992: n_4485 <=  gnd;
delay_3993: a_N456_aNOT_aOUT  <= TRANSPORT a_N456_aNOT_aIN  ;
xor2_3994: a_N456_aNOT_aIN <=  n_4488  XOR n_4497;
or2_3995: n_4488 <=  n_4489  OR n_4493;
and3_3996: n_4489 <=  n_4490  AND n_4491  AND n_4492;
inv_3997: n_4490  <= TRANSPORT NOT a_N1051_aOUT  ;
delay_3998: n_4491  <= TRANSPORT a_N1_aOUT  ;
delay_3999: n_4492  <= TRANSPORT a_N1304_aQ  ;
and3_4000: n_4493 <=  n_4494  AND n_4495  AND n_4496;
inv_4001: n_4494  <= TRANSPORT NOT a_N1050_aOUT  ;
inv_4002: n_4495  <= TRANSPORT NOT a_N1051_aOUT  ;
delay_4003: n_4496  <= TRANSPORT a_N1_aOUT  ;
and1_4004: n_4497 <=  gnd;
delay_4005: a_LC4_A11_aOUT  <= TRANSPORT a_LC4_A11_aIN  ;
xor2_4006: a_LC4_A11_aIN <=  n_4500  XOR n_4509;
or3_4007: n_4500 <=  n_4501  OR n_4503  OR n_4506;
and1_4008: n_4501 <=  n_4502;
inv_4009: n_4502  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and2_4010: n_4503 <=  n_4504  AND n_4505;
inv_4011: n_4504  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
inv_4012: n_4505  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_4013: n_4506 <=  n_4507  AND n_4508;
delay_4014: n_4507  <= TRANSPORT a_N1305_aQ  ;
inv_4015: n_4508  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and1_4016: n_4509 <=  gnd;
delay_4017: a_LC3_A11_aOUT  <= TRANSPORT a_LC3_A11_aIN  ;
xor2_4018: a_LC3_A11_aIN <=  n_4512  XOR n_4521;
or2_4019: n_4512 <=  n_4513  OR n_4517;
and3_4020: n_4513 <=  n_4514  AND n_4515  AND n_4516;
delay_4021: n_4514  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_4022: n_4515  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
delay_4023: n_4516  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and3_4024: n_4517 <=  n_4518  AND n_4519  AND n_4520;
delay_4025: n_4518  <= TRANSPORT a_N1304_aQ  ;
delay_4026: n_4519  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_4027: n_4520  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and1_4028: n_4521 <=  gnd;
delay_4029: a_LC4_A21_aOUT  <= TRANSPORT a_LC4_A21_aIN  ;
xor2_4030: a_LC4_A21_aIN <=  n_4524  XOR n_4534;
or2_4031: n_4524 <=  n_4525  OR n_4529;
and3_4032: n_4525 <=  n_4526  AND n_4527  AND n_4528;
delay_4033: n_4526  <= TRANSPORT a_N1138_aOUT  ;
delay_4034: n_4527  <= TRANSPORT a_N1305_aQ  ;
inv_4035: n_4528  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and3_4036: n_4529 <=  n_4530  AND n_4531  AND n_4533;
delay_4037: n_4530  <= TRANSPORT a_N1138_aOUT  ;
delay_4038: n_4531  <= TRANSPORT a_N1306_aQ  ;
delay_4039: n_4533  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_4040: n_4534 <=  gnd;
delay_4041: a_N1101_aNOT_aOUT  <= TRANSPORT a_N1101_aNOT_aIN  ;
xor2_4042: a_N1101_aNOT_aIN <=  n_4536  XOR n_4545;
or3_4043: n_4536 <=  n_4537  OR n_4540  OR n_4543;
and2_4044: n_4537 <=  n_4538  AND n_4539;
delay_4045: n_4538  <= TRANSPORT a_N456_aNOT_aOUT  ;
delay_4046: n_4539  <= TRANSPORT a_LC4_A11_aOUT  ;
and2_4047: n_4540 <=  n_4541  AND n_4542;
delay_4048: n_4541  <= TRANSPORT a_LC4_A11_aOUT  ;
delay_4049: n_4542  <= TRANSPORT a_LC3_A11_aOUT  ;
and1_4050: n_4543 <=  n_4544;
delay_4051: n_4544  <= TRANSPORT a_LC4_A21_aOUT  ;
and1_4052: n_4545 <=  gnd;
delay_4053: a_N145_aNOT_aOUT  <= TRANSPORT a_N145_aNOT_aIN  ;
xor2_4054: a_N145_aNOT_aIN <=  n_4548  XOR n_4552;
or1_4055: n_4548 <=  n_4549;
and2_4056: n_4549 <=  n_4550  AND n_4551;
inv_4057: n_4550  <= TRANSPORT NOT a_N83_aOUT  ;
delay_4058: n_4551  <= TRANSPORT a_N1101_aNOT_aOUT  ;
and1_4059: n_4552 <=  gnd;
delay_4060: a_N161_aOUT  <= TRANSPORT a_N161_aIN  ;
xor2_4061: a_N161_aIN <=  n_4555  XOR n_4562;
or2_4062: n_4555 <=  n_4556  OR n_4559;
and2_4063: n_4556 <=  n_4557  AND n_4558;
delay_4064: n_4557  <= TRANSPORT a_N1177_aOUT  ;
delay_4065: n_4558  <= TRANSPORT a_N145_aNOT_aOUT  ;
and2_4066: n_4559 <=  n_4560  AND n_4561;
inv_4067: n_4560  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4068: n_4561  <= TRANSPORT a_SRXREG_F1_G_aQ  ;
and1_4069: n_4562 <=  gnd;
delay_4070: a_LC5_A2_aOUT  <= TRANSPORT a_LC5_A2_aIN  ;
xor2_4071: a_LC5_A2_aIN <=  n_4565  XOR n_4574;
or2_4072: n_4565 <=  n_4566  OR n_4570;
and3_4073: n_4566 <=  n_4567  AND n_4568  AND n_4569;
delay_4074: n_4567  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
delay_4075: n_4568  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
inv_4076: n_4569  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and3_4077: n_4570 <=  n_4571  AND n_4572  AND n_4573;
delay_4078: n_4571  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_4079: n_4572  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
delay_4080: n_4573  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_4081: n_4574 <=  gnd;
delay_4082: a_LC1_A21_aOUT  <= TRANSPORT a_LC1_A21_aIN  ;
xor2_4083: a_LC1_A21_aIN <=  n_4577  XOR n_4585;
or2_4084: n_4577 <=  n_4578  OR n_4582;
and2_4085: n_4578 <=  n_4579  AND n_4580;
delay_4086: n_4579  <= TRANSPORT a_N1052_aOUT  ;
delay_4087: n_4580  <= TRANSPORT a_N1307_aQ  ;
and2_4088: n_4582 <=  n_4583  AND n_4584;
delay_4089: n_4583  <= TRANSPORT a_LC5_A2_aOUT  ;
delay_4090: n_4584  <= TRANSPORT a_N1306_aQ  ;
and1_4091: n_4585 <=  gnd;
delay_4092: a_LC5_A21_aOUT  <= TRANSPORT a_LC5_A21_aIN  ;
xor2_4093: a_LC5_A21_aIN <=  n_4588  XOR n_4595;
or2_4094: n_4588 <=  n_4589  OR n_4592;
and2_4095: n_4589 <=  n_4590  AND n_4591;
delay_4096: n_4590  <= TRANSPORT a_N35_aNOT_aOUT  ;
delay_4097: n_4591  <= TRANSPORT a_N1303_aQ  ;
and2_4098: n_4592 <=  n_4593  AND n_4594;
inv_4099: n_4593  <= TRANSPORT NOT a_N35_aNOT_aOUT  ;
delay_4100: n_4594  <= TRANSPORT a_N1304_aQ  ;
and1_4101: n_4595 <=  gnd;
delay_4102: a_LC2_A21_aOUT  <= TRANSPORT a_LC2_A21_aIN  ;
xor2_4103: a_LC2_A21_aIN <=  n_4598  XOR n_4609;
or3_4104: n_4598 <=  n_4599  OR n_4603  OR n_4606;
and3_4105: n_4599 <=  n_4600  AND n_4601  AND n_4602;
inv_4106: n_4600  <= TRANSPORT NOT a_N1050_aOUT  ;
inv_4107: n_4601  <= TRANSPORT NOT a_N1051_aOUT  ;
delay_4108: n_4602  <= TRANSPORT a_LC5_A21_aOUT  ;
and2_4109: n_4603 <=  n_4604  AND n_4605;
delay_4110: n_4604  <= TRANSPORT a_N1051_aOUT  ;
delay_4111: n_4605  <= TRANSPORT a_N1305_aQ  ;
and2_4112: n_4606 <=  n_4607  AND n_4608;
delay_4113: n_4607  <= TRANSPORT a_N1050_aOUT  ;
delay_4114: n_4608  <= TRANSPORT a_N1305_aQ  ;
and1_4115: n_4609 <=  gnd;
delay_4116: a_N1100_aNOT_aOUT  <= TRANSPORT a_N1100_aNOT_aIN  ;
xor2_4117: a_N1100_aNOT_aIN <=  n_4611  XOR n_4618;
or2_4118: n_4611 <=  n_4612  OR n_4614;
and1_4119: n_4612 <=  n_4613;
delay_4120: n_4613  <= TRANSPORT a_LC1_A21_aOUT  ;
and3_4121: n_4614 <=  n_4615  AND n_4616  AND n_4617;
inv_4122: n_4615  <= TRANSPORT NOT a_N1052_aOUT  ;
inv_4123: n_4616  <= TRANSPORT NOT a_N54_aOUT  ;
delay_4124: n_4617  <= TRANSPORT a_LC2_A21_aOUT  ;
and1_4125: n_4618 <=  gnd;
delay_4126: a_N1203_aOUT  <= TRANSPORT a_N1203_aIN  ;
xor2_4127: a_N1203_aIN <=  n_4621  XOR n_4638;
or4_4128: n_4621 <=  n_4622  OR n_4626  OR n_4630  OR n_4634;
and3_4129: n_4622 <=  n_4623  AND n_4624  AND n_4625;
delay_4130: n_4623  <= TRANSPORT a_N676_aOUT  ;
delay_4131: n_4624  <= TRANSPORT a_N1100_aNOT_aOUT  ;
inv_4132: n_4625  <= TRANSPORT NOT a_SSYNC1_F0_G_aQ  ;
and3_4133: n_4626 <=  n_4627  AND n_4628  AND n_4629;
delay_4134: n_4627  <= TRANSPORT a_N676_aOUT  ;
inv_4135: n_4628  <= TRANSPORT NOT a_N1100_aNOT_aOUT  ;
delay_4136: n_4629  <= TRANSPORT a_SSYNC1_F0_G_aQ  ;
and3_4137: n_4630 <=  n_4631  AND n_4632  AND n_4633;
inv_4138: n_4631  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4139: n_4632  <= TRANSPORT NOT a_SSYNC1_F0_G_aQ  ;
delay_4140: n_4633  <= TRANSPORT a_SRXREG_F0_G_aQ  ;
and3_4141: n_4634 <=  n_4635  AND n_4636  AND n_4637;
inv_4142: n_4635  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4143: n_4636  <= TRANSPORT a_SSYNC1_F0_G_aQ  ;
inv_4144: n_4637  <= TRANSPORT NOT a_SRXREG_F0_G_aQ  ;
and1_4145: n_4638 <=  gnd;
delay_4146: a_LC4_B9_aNOT_aOUT  <= TRANSPORT a_LC4_B9_aNOT_aIN  ;
xor2_4147: a_LC4_B9_aNOT_aIN <=  n_4641  XOR n_4652;
or4_4148: n_4641 <=  n_4642  OR n_4644  OR n_4647  OR n_4650;
and1_4149: n_4642 <=  n_4643;
delay_4150: n_4643  <= TRANSPORT a_N1205_aOUT  ;
and2_4151: n_4644 <=  n_4645  AND n_4646;
inv_4152: n_4645  <= TRANSPORT NOT a_SSYNC1_F1_G_aQ  ;
delay_4153: n_4646  <= TRANSPORT a_N161_aOUT  ;
and2_4154: n_4647 <=  n_4648  AND n_4649;
delay_4155: n_4648  <= TRANSPORT a_SSYNC1_F1_G_aQ  ;
inv_4156: n_4649  <= TRANSPORT NOT a_N161_aOUT  ;
and1_4157: n_4650 <=  n_4651;
delay_4158: n_4651  <= TRANSPORT a_N1203_aOUT  ;
and1_4159: n_4652 <=  gnd;
delay_4160: a_LC2_A10_aOUT  <= TRANSPORT a_LC2_A10_aIN  ;
xor2_4161: a_LC2_A10_aIN <=  n_4655  XOR n_4663;
or2_4162: n_4655 <=  n_4656  OR n_4659;
and2_4163: n_4656 <=  n_4657  AND n_4658;
delay_4164: n_4657  <= TRANSPORT a_N1998_aQ  ;
inv_4165: n_4658  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_4166: n_4659 <=  n_4660  AND n_4662;
delay_4167: n_4660  <= TRANSPORT a_N1300_aQ  ;
delay_4168: n_4662  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_4169: n_4663 <=  gnd;
delay_4170: a_N1039_aNOT_aOUT  <= TRANSPORT a_N1039_aNOT_aIN  ;
xor2_4171: a_N1039_aNOT_aIN <=  n_4666  XOR n_4671;
or1_4172: n_4666 <=  n_4667;
and3_4173: n_4667 <=  n_4668  AND n_4669  AND n_4670;
delay_4174: n_4668  <= TRANSPORT a_LC2_A10_aOUT  ;
inv_4175: n_4669  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
delay_4176: n_4670  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_4177: n_4671 <=  gnd;
delay_4178: a_N398_aOUT  <= TRANSPORT a_N398_aIN  ;
xor2_4179: a_N398_aIN <=  n_4674  XOR n_4681;
or3_4180: n_4674 <=  n_4675  OR n_4677  OR n_4679;
and1_4181: n_4675 <=  n_4676;
inv_4182: n_4676  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_4183: n_4677 <=  n_4678;
delay_4184: n_4678  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_4185: n_4679 <=  n_4680;
inv_4186: n_4680  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and1_4187: n_4681 <=  gnd;
delay_4188: a_LC6_A4_aOUT  <= TRANSPORT a_LC6_A4_aIN  ;
xor2_4189: a_LC6_A4_aIN <=  n_4684  XOR n_4697;
or4_4190: n_4684 <=  n_4685  OR n_4688  OR n_4691  OR n_4694;
and2_4191: n_4685 <=  n_4686  AND n_4687;
delay_4192: n_4686  <= TRANSPORT a_N1301_aQ  ;
delay_4193: n_4687  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_4194: n_4688 <=  n_4689  AND n_4690;
inv_4195: n_4689  <= TRANSPORT NOT a_N1138_aOUT  ;
delay_4196: n_4690  <= TRANSPORT a_N1301_aQ  ;
and2_4197: n_4691 <=  n_4692  AND n_4693;
delay_4198: n_4692  <= TRANSPORT a_N398_aOUT  ;
delay_4199: n_4693  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_4200: n_4694 <=  n_4695  AND n_4696;
inv_4201: n_4695  <= TRANSPORT NOT a_N1138_aOUT  ;
delay_4202: n_4696  <= TRANSPORT a_N398_aOUT  ;
and1_4203: n_4697 <=  gnd;
delay_4204: a_N1040_aNOT_aOUT  <= TRANSPORT a_N1040_aNOT_aIN  ;
xor2_4205: a_N1040_aNOT_aIN <=  n_4700  XOR n_4706;
or1_4206: n_4700 <=  n_4701;
and4_4207: n_4701 <=  n_4702  AND n_4703  AND n_4704  AND n_4705;
delay_4208: n_4702  <= TRANSPORT a_N1300_aQ  ;
delay_4209: n_4703  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_4210: n_4704  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
inv_4211: n_4705  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_4212: n_4706 <=  gnd;
delay_4213: a_N687_aNOT_aOUT  <= TRANSPORT a_N687_aNOT_aIN  ;
xor2_4214: a_N687_aNOT_aIN <=  n_4709  XOR n_4719;
or3_4215: n_4709 <=  n_4710  OR n_4713  OR n_4716;
and2_4216: n_4710 <=  n_4711  AND n_4712;
delay_4217: n_4711  <= TRANSPORT a_N1039_aNOT_aOUT  ;
delay_4218: n_4712  <= TRANSPORT a_LC6_A4_aOUT  ;
and2_4219: n_4713 <=  n_4714  AND n_4715;
inv_4220: n_4714  <= TRANSPORT NOT a_N398_aOUT  ;
delay_4221: n_4715  <= TRANSPORT a_LC6_A4_aOUT  ;
and2_4222: n_4716 <=  n_4717  AND n_4718;
delay_4223: n_4717  <= TRANSPORT a_LC6_A4_aOUT  ;
delay_4224: n_4718  <= TRANSPORT a_N1040_aNOT_aOUT  ;
and1_4225: n_4719 <=  gnd;
delay_4226: a_N1041_aNOT_aOUT  <= TRANSPORT a_N1041_aNOT_aIN  ;
xor2_4227: a_N1041_aNOT_aIN <=  n_4722  XOR n_4727;
or1_4228: n_4722 <=  n_4723;
and3_4229: n_4723 <=  n_4724  AND n_4725  AND n_4726;
delay_4230: n_4724  <= TRANSPORT a_N1138_aOUT  ;
delay_4231: n_4725  <= TRANSPORT a_N1301_aQ  ;
inv_4232: n_4726  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_4233: n_4727 <=  gnd;
delay_4234: a_N1105_aNOT_aOUT  <= TRANSPORT a_N1105_aNOT_aIN  ;
xor2_4235: a_N1105_aNOT_aIN <=  n_4729  XOR n_4739;
or3_4236: n_4729 <=  n_4730  OR n_4733  OR n_4736;
and2_4237: n_4730 <=  n_4731  AND n_4732;
inv_4238: n_4731  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4239: n_4732  <= TRANSPORT a_N687_aNOT_aOUT  ;
and2_4240: n_4733 <=  n_4734  AND n_4735;
inv_4241: n_4734  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4242: n_4735  <= TRANSPORT a_N1041_aNOT_aOUT  ;
and2_4243: n_4736 <=  n_4737  AND n_4738;
delay_4244: n_4737  <= TRANSPORT a_N1052_aOUT  ;
delay_4245: n_4738  <= TRANSPORT a_N1302_aQ  ;
and1_4246: n_4739 <=  gnd;
delay_4247: a_N144_aNOT_aOUT  <= TRANSPORT a_N144_aNOT_aIN  ;
xor2_4248: a_N144_aNOT_aIN <=  n_4742  XOR n_4746;
or1_4249: n_4742 <=  n_4743;
and2_4250: n_4743 <=  n_4744  AND n_4745;
inv_4251: n_4744  <= TRANSPORT NOT a_N83_aOUT  ;
delay_4252: n_4745  <= TRANSPORT a_N1105_aNOT_aOUT  ;
and1_4253: n_4746 <=  gnd;
delay_4254: a_N165_aOUT  <= TRANSPORT a_N165_aIN  ;
xor2_4255: a_N165_aIN <=  n_4749  XOR n_4756;
or2_4256: n_4749 <=  n_4750  OR n_4753;
and2_4257: n_4750 <=  n_4751  AND n_4752;
delay_4258: n_4751  <= TRANSPORT a_N1177_aOUT  ;
delay_4259: n_4752  <= TRANSPORT a_N144_aNOT_aOUT  ;
and2_4260: n_4753 <=  n_4754  AND n_4755;
inv_4261: n_4754  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4262: n_4755  <= TRANSPORT a_SRXREG_F5_G_aQ  ;
and1_4263: n_4756 <=  gnd;
delay_4264: a_LC5_C12_aNOT_aOUT  <= TRANSPORT a_LC5_C12_aNOT_aIN  ;
xor2_4265: a_LC5_C12_aNOT_aIN <=  n_4759  XOR n_4772;
or4_4266: n_4759 <=  n_4760  OR n_4762  OR n_4766  OR n_4769;
and1_4267: n_4760 <=  n_4761;
delay_4268: n_4761  <= TRANSPORT a_LC4_B9_aNOT_aOUT  ;
and3_4269: n_4762 <=  n_4763  AND n_4764  AND n_4765;
delay_4270: n_4763  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_4271: n_4764  <= TRANSPORT a_SSYNC1_F5_G_aQ  ;
inv_4272: n_4765  <= TRANSPORT NOT a_N165_aOUT  ;
and2_4273: n_4766 <=  n_4767  AND n_4768;
inv_4274: n_4767  <= TRANSPORT NOT a_SSYNC1_F5_G_aQ  ;
delay_4275: n_4768  <= TRANSPORT a_N165_aOUT  ;
and2_4276: n_4769 <=  n_4770  AND n_4771;
inv_4277: n_4770  <= TRANSPORT NOT a_N1134_aNOT_aOUT  ;
delay_4278: n_4771  <= TRANSPORT a_N165_aOUT  ;
and1_4279: n_4772 <=  gnd;
delay_4280: a_N461_aNOT_aOUT  <= TRANSPORT a_N461_aNOT_aIN  ;
xor2_4281: a_N461_aNOT_aIN <=  n_4775  XOR n_4786;
or3_4282: n_4775 <=  n_4776  OR n_4780  OR n_4783;
and3_4283: n_4776 <=  n_4777  AND n_4778  AND n_4779;
inv_4284: n_4777  <= TRANSPORT NOT a_N1134_aNOT_aOUT  ;
delay_4285: n_4778  <= TRANSPORT a_N1301_aQ  ;
delay_4286: n_4779  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_4287: n_4780 <=  n_4781  AND n_4782;
delay_4288: n_4781  <= TRANSPORT a_N1300_aQ  ;
inv_4289: n_4782  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_4290: n_4783 <=  n_4784  AND n_4785;
delay_4291: n_4784  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_4292: n_4785  <= TRANSPORT a_N1300_aQ  ;
and1_4293: n_4786 <=  gnd;
delay_4294: a_N458_aNOT_aOUT  <= TRANSPORT a_N458_aNOT_aIN  ;
xor2_4295: a_N458_aNOT_aIN <=  n_4789  XOR n_4793;
or1_4296: n_4789 <=  n_4790;
and2_4297: n_4790 <=  n_4791  AND n_4792;
delay_4298: n_4791  <= TRANSPORT a_N1049_aNOT_aOUT  ;
delay_4299: n_4792  <= TRANSPORT a_N461_aNOT_aOUT  ;
and1_4300: n_4793 <=  gnd;
delay_4301: a_N22_aNOT_aOUT  <= TRANSPORT a_N22_aNOT_aIN  ;
xor2_4302: a_N22_aNOT_aIN <=  n_4796  XOR n_4801;
or1_4303: n_4796 <=  n_4797;
and3_4304: n_4797 <=  n_4798  AND n_4799  AND n_4800;
delay_4305: n_4798  <= TRANSPORT a_N1301_aQ  ;
inv_4306: n_4799  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
delay_4307: n_4800  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_4308: n_4801 <=  gnd;
delay_4309: a_N20_aNOT_aOUT  <= TRANSPORT a_N20_aNOT_aIN  ;
xor2_4310: a_N20_aNOT_aIN <=  n_4804  XOR n_4813;
or2_4311: n_4804 <=  n_4805  OR n_4809;
and3_4312: n_4805 <=  n_4806  AND n_4807  AND n_4808;
inv_4313: n_4806  <= TRANSPORT NOT a_N1050_aOUT  ;
inv_4314: n_4807  <= TRANSPORT NOT a_N1051_aOUT  ;
delay_4315: n_4808  <= TRANSPORT a_N458_aNOT_aOUT  ;
and3_4316: n_4809 <=  n_4810  AND n_4811  AND n_4812;
inv_4317: n_4810  <= TRANSPORT NOT a_N1050_aOUT  ;
inv_4318: n_4811  <= TRANSPORT NOT a_N1051_aOUT  ;
delay_4319: n_4812  <= TRANSPORT a_N22_aNOT_aOUT  ;
and1_4320: n_4813 <=  gnd;
delay_4321: a_N19_aNOT_aOUT  <= TRANSPORT a_N19_aNOT_aIN  ;
xor2_4322: a_N19_aNOT_aIN <=  n_4816  XOR n_4823;
or2_4323: n_4816 <=  n_4817  OR n_4820;
and2_4324: n_4817 <=  n_4818  AND n_4819;
delay_4325: n_4818  <= TRANSPORT a_N1051_aOUT  ;
delay_4326: n_4819  <= TRANSPORT a_N1302_aQ  ;
and2_4327: n_4820 <=  n_4821  AND n_4822;
delay_4328: n_4821  <= TRANSPORT a_N1050_aOUT  ;
delay_4329: n_4822  <= TRANSPORT a_N1302_aQ  ;
and1_4330: n_4823 <=  gnd;
delay_4331: a_N55_aNOT_aOUT  <= TRANSPORT a_N55_aNOT_aIN  ;
xor2_4332: a_N55_aNOT_aIN <=  n_4826  XOR n_4833;
or2_4333: n_4826 <=  n_4827  OR n_4830;
and2_4334: n_4827 <=  n_4828  AND n_4829;
inv_4335: n_4828  <= TRANSPORT NOT a_N54_aOUT  ;
delay_4336: n_4829  <= TRANSPORT a_N20_aNOT_aOUT  ;
and2_4337: n_4830 <=  n_4831  AND n_4832;
inv_4338: n_4831  <= TRANSPORT NOT a_N54_aOUT  ;
delay_4339: n_4832  <= TRANSPORT a_N19_aNOT_aOUT  ;
and1_4340: n_4833 <=  gnd;
delay_4341: a_N56_aNOT_aOUT  <= TRANSPORT a_N56_aNOT_aIN  ;
xor2_4342: a_N56_aNOT_aIN <=  n_4836  XOR n_4840;
or1_4343: n_4836 <=  n_4837;
and2_4344: n_4837 <=  n_4838  AND n_4839;
delay_4345: n_4838  <= TRANSPORT a_N54_aOUT  ;
delay_4346: n_4839  <= TRANSPORT a_N1303_aQ  ;
and1_4347: n_4840 <=  gnd;
delay_4348: a_N1103_aNOT_aOUT  <= TRANSPORT a_N1103_aNOT_aIN  ;
xor2_4349: a_N1103_aNOT_aIN <=  n_4842  XOR n_4852;
or3_4350: n_4842 <=  n_4843  OR n_4846  OR n_4849;
and2_4351: n_4843 <=  n_4844  AND n_4845;
inv_4352: n_4844  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4353: n_4845  <= TRANSPORT a_N55_aNOT_aOUT  ;
and2_4354: n_4846 <=  n_4847  AND n_4848;
inv_4355: n_4847  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4356: n_4848  <= TRANSPORT a_N56_aNOT_aOUT  ;
and2_4357: n_4849 <=  n_4850  AND n_4851;
delay_4358: n_4850  <= TRANSPORT a_N1052_aOUT  ;
delay_4359: n_4851  <= TRANSPORT a_N1304_aQ  ;
and1_4360: n_4852 <=  gnd;
delay_4361: a_N1206_aOUT  <= TRANSPORT a_N1206_aIN  ;
xor2_4362: a_N1206_aIN <=  n_4855  XOR n_4872;
or4_4363: n_4855 <=  n_4856  OR n_4860  OR n_4864  OR n_4868;
and3_4364: n_4856 <=  n_4857  AND n_4858  AND n_4859;
inv_4365: n_4857  <= TRANSPORT NOT a_SSYNC1_F3_G_aQ  ;
delay_4366: n_4858  <= TRANSPORT a_N676_aOUT  ;
delay_4367: n_4859  <= TRANSPORT a_N1103_aNOT_aOUT  ;
and3_4368: n_4860 <=  n_4861  AND n_4862  AND n_4863;
inv_4369: n_4861  <= TRANSPORT NOT a_SSYNC1_F3_G_aQ  ;
inv_4370: n_4862  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4371: n_4863  <= TRANSPORT a_SRXREG_F3_G_aQ  ;
and3_4372: n_4864 <=  n_4865  AND n_4866  AND n_4867;
delay_4373: n_4865  <= TRANSPORT a_SSYNC1_F3_G_aQ  ;
delay_4374: n_4866  <= TRANSPORT a_N676_aOUT  ;
inv_4375: n_4867  <= TRANSPORT NOT a_N1103_aNOT_aOUT  ;
and3_4376: n_4868 <=  n_4869  AND n_4870  AND n_4871;
delay_4377: n_4869  <= TRANSPORT a_SSYNC1_F3_G_aQ  ;
inv_4378: n_4870  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4379: n_4871  <= TRANSPORT NOT a_SRXREG_F3_G_aQ  ;
and1_4380: n_4872 <=  gnd;
delay_4381: a_N96_aOUT  <= TRANSPORT a_N96_aIN  ;
xor2_4382: a_N96_aIN <=  n_4874  XOR n_4879;
or1_4383: n_4874 <=  n_4875;
and3_4384: n_4875 <=  n_4876  AND n_4877  AND n_4878;
delay_4385: n_4876  <= TRANSPORT a_LC2_A10_aOUT  ;
delay_4386: n_4877  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
delay_4387: n_4878  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_4388: n_4879 <=  gnd;
delay_4389: a_N166_aOUT  <= TRANSPORT a_N166_aIN  ;
xor2_4390: a_N166_aIN <=  n_4882  XOR n_4889;
or2_4391: n_4882 <=  n_4883  OR n_4886;
and2_4392: n_4883 <=  n_4884  AND n_4885;
delay_4393: n_4884  <= TRANSPORT a_N676_aOUT  ;
delay_4394: n_4885  <= TRANSPORT a_N96_aOUT  ;
and2_4395: n_4886 <=  n_4887  AND n_4888;
inv_4396: n_4887  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4397: n_4888  <= TRANSPORT a_SRXREG_F7_G_aQ  ;
and1_4398: n_4889 <=  gnd;
delay_4399: a_LC2_C11_aNOT_aOUT  <= TRANSPORT a_LC2_C11_aNOT_aIN  ;
xor2_4400: a_LC2_C11_aNOT_aIN <=  n_4892  XOR n_4905;
or4_4401: n_4892 <=  n_4893  OR n_4895  OR n_4899  OR n_4902;
and1_4402: n_4893 <=  n_4894;
delay_4403: n_4894  <= TRANSPORT a_N1206_aOUT  ;
and3_4404: n_4895 <=  n_4896  AND n_4897  AND n_4898;
delay_4405: n_4896  <= TRANSPORT a_N1138_aOUT  ;
delay_4406: n_4897  <= TRANSPORT a_SSYNC1_F7_G_aQ  ;
inv_4407: n_4898  <= TRANSPORT NOT a_N166_aOUT  ;
and2_4408: n_4899 <=  n_4900  AND n_4901;
inv_4409: n_4900  <= TRANSPORT NOT a_SSYNC1_F7_G_aQ  ;
delay_4410: n_4901  <= TRANSPORT a_N166_aOUT  ;
and2_4411: n_4902 <=  n_4903  AND n_4904;
inv_4412: n_4903  <= TRANSPORT NOT a_N1138_aOUT  ;
delay_4413: n_4904  <= TRANSPORT a_N166_aOUT  ;
and1_4414: n_4905 <=  gnd;
delay_4415: a_LC3_A19_aOUT  <= TRANSPORT a_LC3_A19_aIN  ;
xor2_4416: a_LC3_A19_aIN <=  n_4908  XOR n_4913;
or1_4417: n_4908 <=  n_4909;
and3_4418: n_4909 <=  n_4910  AND n_4911  AND n_4912;
delay_4419: n_4910  <= TRANSPORT a_N1138_aOUT  ;
delay_4420: n_4911  <= TRANSPORT a_N1300_aQ  ;
inv_4421: n_4912  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_4422: n_4913 <=  gnd;
delay_4423: a_LC1_A19_aOUT  <= TRANSPORT a_LC1_A19_aIN  ;
xor2_4424: a_LC1_A19_aIN <=  n_4916  XOR n_4921;
or1_4425: n_4916 <=  n_4917;
and3_4426: n_4917 <=  n_4918  AND n_4919  AND n_4920;
delay_4427: n_4918  <= TRANSPORT a_LC2_A10_aOUT  ;
delay_4428: n_4919  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
inv_4429: n_4920  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and1_4430: n_4921 <=  gnd;
delay_4431: a_N1106_aNOT_aOUT  <= TRANSPORT a_N1106_aNOT_aIN  ;
xor2_4432: a_N1106_aNOT_aIN <=  n_4923  XOR n_4933;
or3_4433: n_4923 <=  n_4924  OR n_4927  OR n_4930;
and2_4434: n_4924 <=  n_4925  AND n_4926;
delay_4435: n_4925  <= TRANSPORT a_N1052_aOUT  ;
delay_4436: n_4926  <= TRANSPORT a_N1301_aQ  ;
and2_4437: n_4927 <=  n_4928  AND n_4929;
inv_4438: n_4928  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4439: n_4929  <= TRANSPORT a_LC3_A19_aOUT  ;
and2_4440: n_4930 <=  n_4931  AND n_4932;
inv_4441: n_4931  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4442: n_4932  <= TRANSPORT a_LC1_A19_aOUT  ;
and1_4443: n_4933 <=  gnd;
delay_4444: a_N686_aOUT  <= TRANSPORT a_N686_aIN  ;
xor2_4445: a_N686_aIN <=  n_4936  XOR n_4943;
or2_4446: n_4936 <=  n_4937  OR n_4940;
and2_4447: n_4937 <=  n_4938  AND n_4939;
delay_4448: n_4938  <= TRANSPORT a_N676_aOUT  ;
delay_4449: n_4939  <= TRANSPORT a_N1106_aNOT_aOUT  ;
and2_4450: n_4940 <=  n_4941  AND n_4942;
inv_4451: n_4941  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4452: n_4942  <= TRANSPORT a_SRXREG_F6_G_aQ  ;
and1_4453: n_4943 <=  gnd;
delay_4454: a_N1077_aOUT  <= TRANSPORT a_N1077_aIN  ;
xor2_4455: a_N1077_aIN <=  n_4946  XOR n_4957;
or3_4456: n_4946 <=  n_4947  OR n_4951  OR n_4954;
and3_4457: n_4947 <=  n_4948  AND n_4949  AND n_4950;
delay_4458: n_4948  <= TRANSPORT a_SSYNC1_F6_G_aQ  ;
inv_4459: n_4949  <= TRANSPORT NOT a_N686_aOUT  ;
delay_4460: n_4950  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and2_4461: n_4951 <=  n_4952  AND n_4953;
delay_4462: n_4952  <= TRANSPORT a_N686_aOUT  ;
inv_4463: n_4953  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and2_4464: n_4954 <=  n_4955  AND n_4956;
inv_4465: n_4955  <= TRANSPORT NOT a_SSYNC1_F6_G_aQ  ;
delay_4466: n_4956  <= TRANSPORT a_N686_aOUT  ;
and1_4467: n_4957 <=  gnd;
delay_4468: a_N694_aNOT_aOUT  <= TRANSPORT a_N694_aNOT_aIN  ;
xor2_4469: a_N694_aNOT_aIN <=  n_4960  XOR n_4967;
or2_4470: n_4960 <=  n_4961  OR n_4964;
and2_4471: n_4961 <=  n_4962  AND n_4963;
delay_4472: n_4962  <= TRANSPORT a_N1051_aOUT  ;
delay_4473: n_4963  <= TRANSPORT a_N1301_aQ  ;
and2_4474: n_4964 <=  n_4965  AND n_4966;
delay_4475: n_4965  <= TRANSPORT a_LC5_A2_aOUT  ;
delay_4476: n_4966  <= TRANSPORT a_N1302_aQ  ;
and1_4477: n_4967 <=  gnd;
delay_4478: a_N696_aNOT_aOUT  <= TRANSPORT a_N696_aNOT_aIN  ;
xor2_4479: a_N696_aNOT_aIN <=  n_4970  XOR n_4977;
or2_4480: n_4970 <=  n_4971  OR n_4974;
and2_4481: n_4971 <=  n_4972  AND n_4973;
delay_4482: n_4972  <= TRANSPORT a_N1300_aQ  ;
inv_4483: n_4973  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_4484: n_4974 <=  n_4975  AND n_4976;
delay_4485: n_4975  <= TRANSPORT a_N1301_aQ  ;
delay_4486: n_4976  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_4487: n_4977 <=  gnd;
delay_4488: a_LC6_A19_aOUT  <= TRANSPORT a_LC6_A19_aIN  ;
xor2_4489: a_LC6_A19_aIN <=  n_4980  XOR n_4989;
or2_4490: n_4980 <=  n_4981  OR n_4985;
and3_4491: n_4981 <=  n_4982  AND n_4983  AND n_4984;
delay_4492: n_4982  <= TRANSPORT a_LC2_A10_aOUT  ;
inv_4493: n_4983  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
inv_4494: n_4984  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
and3_4495: n_4985 <=  n_4986  AND n_4987  AND n_4988;
delay_4496: n_4986  <= TRANSPORT a_N696_aNOT_aOUT  ;
inv_4497: n_4987  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
delay_4498: n_4988  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
and1_4499: n_4989 <=  gnd;
delay_4500: a_N1104_aNOT_aOUT  <= TRANSPORT a_N1104_aNOT_aIN  ;
xor2_4501: a_N1104_aNOT_aIN <=  n_4991  XOR n_5000;
or3_4502: n_4991 <=  n_4992  OR n_4995  OR n_4998;
and2_4503: n_4992 <=  n_4993  AND n_4994;
inv_4504: n_4993  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_4505: n_4994  <= TRANSPORT a_N694_aNOT_aOUT  ;
and2_4506: n_4995 <=  n_4996  AND n_4997;
delay_4507: n_4996  <= TRANSPORT a_N1052_aOUT  ;
delay_4508: n_4997  <= TRANSPORT a_N1303_aQ  ;
and1_4509: n_4998 <=  n_4999;
delay_4510: n_4999  <= TRANSPORT a_LC6_A19_aOUT  ;
and1_4511: n_5000 <=  gnd;
delay_4512: a_N1207_aOUT  <= TRANSPORT a_N1207_aIN  ;
xor2_4513: a_N1207_aIN <=  n_5003  XOR n_5020;
or4_4514: n_5003 <=  n_5004  OR n_5008  OR n_5012  OR n_5016;
and3_4515: n_5004 <=  n_5005  AND n_5006  AND n_5007;
inv_4516: n_5005  <= TRANSPORT NOT a_SSYNC1_F4_G_aQ  ;
delay_4517: n_5006  <= TRANSPORT a_N676_aOUT  ;
delay_4518: n_5007  <= TRANSPORT a_N1104_aNOT_aOUT  ;
and3_4519: n_5008 <=  n_5009  AND n_5010  AND n_5011;
inv_4520: n_5009  <= TRANSPORT NOT a_SSYNC1_F4_G_aQ  ;
inv_4521: n_5010  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4522: n_5011  <= TRANSPORT a_SRXREG_F4_G_aQ  ;
and3_4523: n_5012 <=  n_5013  AND n_5014  AND n_5015;
delay_4524: n_5013  <= TRANSPORT a_SSYNC1_F4_G_aQ  ;
inv_4525: n_5014  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4526: n_5015  <= TRANSPORT NOT a_SRXREG_F4_G_aQ  ;
and3_4527: n_5016 <=  n_5017  AND n_5018  AND n_5019;
delay_4528: n_5017  <= TRANSPORT a_SSYNC1_F4_G_aQ  ;
delay_4529: n_5018  <= TRANSPORT a_N676_aOUT  ;
inv_4530: n_5019  <= TRANSPORT NOT a_N1104_aNOT_aOUT  ;
and1_4531: n_5020 <=  gnd;
delay_4532: a_N135_aOUT  <= TRANSPORT a_N135_aIN  ;
xor2_4533: a_N135_aIN <=  n_5023  XOR n_5032;
or4_4534: n_5023 <=  n_5024  OR n_5026  OR n_5028  OR n_5030;
and1_4535: n_5024 <=  n_5025;
delay_4536: n_5025  <= TRANSPORT a_LC5_C12_aNOT_aOUT  ;
and1_4537: n_5026 <=  n_5027;
delay_4538: n_5027  <= TRANSPORT a_LC2_C11_aNOT_aOUT  ;
and1_4539: n_5028 <=  n_5029;
delay_4540: n_5029  <= TRANSPORT a_N1077_aOUT  ;
and1_4541: n_5030 <=  n_5031;
delay_4542: n_5031  <= TRANSPORT a_N1207_aOUT  ;
and1_4543: n_5032 <=  gnd;
delay_4544: a_N1038_aNOT_aOUT  <= TRANSPORT a_N1038_aNOT_aIN  ;
xor2_4545: a_N1038_aNOT_aIN <=  n_5035  XOR n_5042;
or3_4546: n_5035 <=  n_5036  OR n_5038  OR n_5040;
and1_4547: n_5036 <=  n_5037;
delay_4548: n_5037  <= TRANSPORT a_N1555_aQ  ;
and1_4549: n_5038 <=  n_5039;
inv_4550: n_5039  <= TRANSPORT NOT a_N1556_aQ  ;
and1_4551: n_5040 <=  n_5041;
delay_4552: n_5041  <= TRANSPORT a_N135_aOUT  ;
and1_4553: n_5042 <=  gnd;
delay_4554: a_N1212_aOUT  <= TRANSPORT a_N1212_aIN  ;
xor2_4555: a_N1212_aIN <=  n_5045  XOR n_5062;
or4_4556: n_5045 <=  n_5046  OR n_5050  OR n_5054  OR n_5058;
and3_4557: n_5046 <=  n_5047  AND n_5048  AND n_5049;
inv_4558: n_5047  <= TRANSPORT NOT a_SSYNC2_F2_G_aQ  ;
delay_4559: n_5048  <= TRANSPORT a_N676_aOUT  ;
delay_4560: n_5049  <= TRANSPORT a_N1102_aNOT_aOUT  ;
and3_4561: n_5050 <=  n_5051  AND n_5052  AND n_5053;
inv_4562: n_5051  <= TRANSPORT NOT a_SSYNC2_F2_G_aQ  ;
inv_4563: n_5052  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4564: n_5053  <= TRANSPORT a_SRXREG_F2_G_aQ  ;
and3_4565: n_5054 <=  n_5055  AND n_5056  AND n_5057;
delay_4566: n_5055  <= TRANSPORT a_SSYNC2_F2_G_aQ  ;
delay_4567: n_5056  <= TRANSPORT a_N676_aOUT  ;
inv_4568: n_5057  <= TRANSPORT NOT a_N1102_aNOT_aOUT  ;
and3_4569: n_5058 <=  n_5059  AND n_5060  AND n_5061;
delay_4570: n_5059  <= TRANSPORT a_SSYNC2_F2_G_aQ  ;
inv_4571: n_5060  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4572: n_5061  <= TRANSPORT NOT a_SRXREG_F2_G_aQ  ;
and1_4573: n_5062 <=  gnd;
delay_4574: a_N1210_aOUT  <= TRANSPORT a_N1210_aIN  ;
xor2_4575: a_N1210_aIN <=  n_5065  XOR n_5082;
or4_4576: n_5065 <=  n_5066  OR n_5070  OR n_5074  OR n_5078;
and3_4577: n_5066 <=  n_5067  AND n_5068  AND n_5069;
delay_4578: n_5067  <= TRANSPORT a_N676_aOUT  ;
delay_4579: n_5068  <= TRANSPORT a_N1100_aNOT_aOUT  ;
inv_4580: n_5069  <= TRANSPORT NOT a_SSYNC2_F0_G_aQ  ;
and3_4581: n_5070 <=  n_5071  AND n_5072  AND n_5073;
delay_4582: n_5071  <= TRANSPORT a_N676_aOUT  ;
inv_4583: n_5072  <= TRANSPORT NOT a_N1100_aNOT_aOUT  ;
delay_4584: n_5073  <= TRANSPORT a_SSYNC2_F0_G_aQ  ;
and3_4585: n_5074 <=  n_5075  AND n_5076  AND n_5077;
inv_4586: n_5075  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4587: n_5076  <= TRANSPORT NOT a_SSYNC2_F0_G_aQ  ;
delay_4588: n_5077  <= TRANSPORT a_SRXREG_F0_G_aQ  ;
and3_4589: n_5078 <=  n_5079  AND n_5080  AND n_5081;
inv_4590: n_5079  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4591: n_5080  <= TRANSPORT a_SSYNC2_F0_G_aQ  ;
inv_4592: n_5081  <= TRANSPORT NOT a_SRXREG_F0_G_aQ  ;
and1_4593: n_5082 <=  gnd;
delay_4594: a_LC2_B9_aOUT  <= TRANSPORT a_LC2_B9_aIN  ;
xor2_4595: a_LC2_B9_aIN <=  n_5085  XOR n_5096;
or4_4596: n_5085 <=  n_5086  OR n_5088  OR n_5091  OR n_5094;
and1_4597: n_5086 <=  n_5087;
delay_4598: n_5087  <= TRANSPORT a_N1212_aOUT  ;
and2_4599: n_5088 <=  n_5089  AND n_5090;
inv_4600: n_5089  <= TRANSPORT NOT a_SSYNC2_F1_G_aQ  ;
delay_4601: n_5090  <= TRANSPORT a_N161_aOUT  ;
and2_4602: n_5091 <=  n_5092  AND n_5093;
delay_4603: n_5092  <= TRANSPORT a_SSYNC2_F1_G_aQ  ;
inv_4604: n_5093  <= TRANSPORT NOT a_N161_aOUT  ;
and1_4605: n_5094 <=  n_5095;
delay_4606: n_5095  <= TRANSPORT a_N1210_aOUT  ;
and1_4607: n_5096 <=  gnd;
delay_4608: a_LC1_C12_aOUT  <= TRANSPORT a_LC1_C12_aIN  ;
xor2_4609: a_LC1_C12_aIN <=  n_5099  XOR n_5112;
or4_4610: n_5099 <=  n_5100  OR n_5102  OR n_5106  OR n_5109;
and1_4611: n_5100 <=  n_5101;
delay_4612: n_5101  <= TRANSPORT a_LC2_B9_aOUT  ;
and3_4613: n_5102 <=  n_5103  AND n_5104  AND n_5105;
delay_4614: n_5103  <= TRANSPORT a_SSYNC2_F6_G_aQ  ;
inv_4615: n_5104  <= TRANSPORT NOT a_N686_aOUT  ;
delay_4616: n_5105  <= TRANSPORT a_SMODE_OUT_F3_G_aQ  ;
and2_4617: n_5106 <=  n_5107  AND n_5108;
delay_4618: n_5107  <= TRANSPORT a_N686_aOUT  ;
inv_4619: n_5108  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and2_4620: n_5109 <=  n_5110  AND n_5111;
inv_4621: n_5110  <= TRANSPORT NOT a_SSYNC2_F6_G_aQ  ;
delay_4622: n_5111  <= TRANSPORT a_N686_aOUT  ;
and1_4623: n_5112 <=  gnd;
delay_4624: a_N1213_aOUT  <= TRANSPORT a_N1213_aIN  ;
xor2_4625: a_N1213_aIN <=  n_5115  XOR n_5132;
or4_4626: n_5115 <=  n_5116  OR n_5120  OR n_5124  OR n_5128;
and3_4627: n_5116 <=  n_5117  AND n_5118  AND n_5119;
inv_4628: n_5117  <= TRANSPORT NOT a_SSYNC2_F3_G_aQ  ;
delay_4629: n_5118  <= TRANSPORT a_N676_aOUT  ;
delay_4630: n_5119  <= TRANSPORT a_N1103_aNOT_aOUT  ;
and3_4631: n_5120 <=  n_5121  AND n_5122  AND n_5123;
inv_4632: n_5121  <= TRANSPORT NOT a_SSYNC2_F3_G_aQ  ;
inv_4633: n_5122  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4634: n_5123  <= TRANSPORT a_SRXREG_F3_G_aQ  ;
and3_4635: n_5124 <=  n_5125  AND n_5126  AND n_5127;
delay_4636: n_5125  <= TRANSPORT a_SSYNC2_F3_G_aQ  ;
delay_4637: n_5126  <= TRANSPORT a_N676_aOUT  ;
inv_4638: n_5127  <= TRANSPORT NOT a_N1103_aNOT_aOUT  ;
and3_4639: n_5128 <=  n_5129  AND n_5130  AND n_5131;
delay_4640: n_5129  <= TRANSPORT a_SSYNC2_F3_G_aQ  ;
inv_4641: n_5130  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4642: n_5131  <= TRANSPORT NOT a_SRXREG_F3_G_aQ  ;
and1_4643: n_5132 <=  gnd;
delay_4644: a_LC1_C11_aOUT  <= TRANSPORT a_LC1_C11_aIN  ;
xor2_4645: a_LC1_C11_aIN <=  n_5135  XOR n_5148;
or4_4646: n_5135 <=  n_5136  OR n_5138  OR n_5142  OR n_5145;
and1_4647: n_5136 <=  n_5137;
delay_4648: n_5137  <= TRANSPORT a_N1213_aOUT  ;
and3_4649: n_5138 <=  n_5139  AND n_5140  AND n_5141;
delay_4650: n_5139  <= TRANSPORT a_N1138_aOUT  ;
delay_4651: n_5140  <= TRANSPORT a_SSYNC2_F7_G_aQ  ;
inv_4652: n_5141  <= TRANSPORT NOT a_N166_aOUT  ;
and2_4653: n_5142 <=  n_5143  AND n_5144;
inv_4654: n_5143  <= TRANSPORT NOT a_SSYNC2_F7_G_aQ  ;
delay_4655: n_5144  <= TRANSPORT a_N166_aOUT  ;
and2_4656: n_5145 <=  n_5146  AND n_5147;
inv_4657: n_5146  <= TRANSPORT NOT a_N1138_aOUT  ;
delay_4658: n_5147  <= TRANSPORT a_N166_aOUT  ;
and1_4659: n_5148 <=  gnd;
delay_4660: a_N1215_aOUT  <= TRANSPORT a_N1215_aIN  ;
xor2_4661: a_N1215_aIN <=  n_5151  XOR n_5162;
or3_4662: n_5151 <=  n_5152  OR n_5156  OR n_5159;
and3_4663: n_5152 <=  n_5153  AND n_5154  AND n_5155;
delay_4664: n_5153  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_4665: n_5154  <= TRANSPORT a_SSYNC2_F5_G_aQ  ;
inv_4666: n_5155  <= TRANSPORT NOT a_N165_aOUT  ;
and2_4667: n_5156 <=  n_5157  AND n_5158;
inv_4668: n_5157  <= TRANSPORT NOT a_SSYNC2_F5_G_aQ  ;
delay_4669: n_5158  <= TRANSPORT a_N165_aOUT  ;
and2_4670: n_5159 <=  n_5160  AND n_5161;
inv_4671: n_5160  <= TRANSPORT NOT a_N1134_aNOT_aOUT  ;
delay_4672: n_5161  <= TRANSPORT a_N165_aOUT  ;
and1_4673: n_5162 <=  gnd;
delay_4674: a_N1214_aOUT  <= TRANSPORT a_N1214_aIN  ;
xor2_4675: a_N1214_aIN <=  n_5165  XOR n_5182;
or4_4676: n_5165 <=  n_5166  OR n_5170  OR n_5174  OR n_5178;
and3_4677: n_5166 <=  n_5167  AND n_5168  AND n_5169;
inv_4678: n_5167  <= TRANSPORT NOT a_SSYNC2_F4_G_aQ  ;
delay_4679: n_5168  <= TRANSPORT a_N676_aOUT  ;
delay_4680: n_5169  <= TRANSPORT a_N1104_aNOT_aOUT  ;
and3_4681: n_5170 <=  n_5171  AND n_5172  AND n_5173;
inv_4682: n_5171  <= TRANSPORT NOT a_SSYNC2_F4_G_aQ  ;
inv_4683: n_5172  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4684: n_5173  <= TRANSPORT a_SRXREG_F4_G_aQ  ;
and3_4685: n_5174 <=  n_5175  AND n_5176  AND n_5177;
delay_4686: n_5175  <= TRANSPORT a_SSYNC2_F4_G_aQ  ;
inv_4687: n_5176  <= TRANSPORT NOT a_N676_aOUT  ;
inv_4688: n_5177  <= TRANSPORT NOT a_SRXREG_F4_G_aQ  ;
and3_4689: n_5178 <=  n_5179  AND n_5180  AND n_5181;
delay_4690: n_5179  <= TRANSPORT a_SSYNC2_F4_G_aQ  ;
delay_4691: n_5180  <= TRANSPORT a_N676_aOUT  ;
inv_4692: n_5181  <= TRANSPORT NOT a_N1104_aNOT_aOUT  ;
and1_4693: n_5182 <=  gnd;
delay_4694: a_N1194_aNOT_aOUT  <= TRANSPORT a_N1194_aNOT_aIN  ;
xor2_4695: a_N1194_aNOT_aIN <=  n_5185  XOR n_5194;
or4_4696: n_5185 <=  n_5186  OR n_5188  OR n_5190  OR n_5192;
and1_4697: n_5186 <=  n_5187;
delay_4698: n_5187  <= TRANSPORT a_LC1_C12_aOUT  ;
and1_4699: n_5188 <=  n_5189;
delay_4700: n_5189  <= TRANSPORT a_LC1_C11_aOUT  ;
and1_4701: n_5190 <=  n_5191;
delay_4702: n_5191  <= TRANSPORT a_N1215_aOUT  ;
and1_4703: n_5192 <=  n_5193;
delay_4704: n_5193  <= TRANSPORT a_N1214_aOUT  ;
and1_4705: n_5194 <=  gnd;
delay_4706: a_N1037_aNOT_aOUT  <= TRANSPORT a_N1037_aNOT_aIN  ;
xor2_4707: a_N1037_aNOT_aIN <=  n_5197  XOR n_5206;
or4_4708: n_5197 <=  n_5198  OR n_5200  OR n_5202  OR n_5204;
and1_4709: n_5198 <=  n_5199;
delay_4710: n_5199  <= TRANSPORT a_N1194_aNOT_aOUT  ;
and1_4711: n_5200 <=  n_5201;
inv_4712: n_5201  <= TRANSPORT NOT a_N1555_aQ  ;
and1_4713: n_5202 <=  n_5203;
delay_4714: n_5203  <= TRANSPORT a_N1556_aQ  ;
and1_4715: n_5204 <=  n_5205;
delay_4716: n_5205  <= TRANSPORT a_N132_aOUT  ;
and1_4717: n_5206 <=  gnd;
delay_4718: a_LC6_A15_aOUT  <= TRANSPORT a_LC6_A15_aIN  ;
xor2_4719: a_LC6_A15_aIN <=  n_5209  XOR n_5217;
or2_4720: n_5209 <=  n_5210  OR n_5214;
and3_4721: n_5210 <=  n_5211  AND n_5212  AND n_5213;
delay_4722: n_5211  <= TRANSPORT a_N1038_aNOT_aOUT  ;
delay_4723: n_5212  <= TRANSPORT a_N1037_aNOT_aOUT  ;
delay_4724: n_5213  <= TRANSPORT nRESET  ;
and2_4725: n_5214 <=  n_5215  AND n_5216;
inv_4726: n_5215  <= TRANSPORT NOT a_N676_aOUT  ;
delay_4727: n_5216  <= TRANSPORT nRESET  ;
and1_4728: n_5217 <=  gnd;
delay_4729: a_N1125_aOUT  <= TRANSPORT a_N1125_aIN  ;
xor2_4730: a_N1125_aIN <=  n_5220  XOR n_5230;
or3_4731: n_5220 <=  n_5221  OR n_5224  OR n_5227;
and2_4732: n_5221 <=  n_5222  AND n_5223;
delay_4733: n_5222  <= TRANSPORT a_N167_aOUT  ;
delay_4734: n_5223  <= TRANSPORT a_LC6_A15_aOUT  ;
and2_4735: n_5224 <=  n_5225  AND n_5226;
delay_4736: n_5225  <= TRANSPORT a_N676_aOUT  ;
delay_4737: n_5226  <= TRANSPORT a_LC6_A15_aOUT  ;
and2_4738: n_5227 <=  n_5228  AND n_5229;
delay_4739: n_5228  <= TRANSPORT a_N83_aOUT  ;
delay_4740: n_5229  <= TRANSPORT a_LC6_A15_aOUT  ;
and1_4741: n_5230 <=  gnd;
delay_4742: a_N86_aOUT  <= TRANSPORT a_N86_aIN  ;
xor2_4743: a_N86_aIN <=  n_5233  XOR n_5239;
or1_4744: n_5233 <=  n_5234;
and4_4745: n_5234 <=  n_5235  AND n_5236  AND n_5237  AND n_5238;
delay_4746: n_5235  <= TRANSPORT a_N127_aOUT  ;
delay_4747: n_5236  <= TRANSPORT a_N59_aQ  ;
inv_4748: n_5237  <= TRANSPORT NOT a_N62_aQ  ;
inv_4749: n_5238  <= TRANSPORT NOT a_N63_aQ  ;
and1_4750: n_5239 <=  gnd;
delay_4751: a_N91_aOUT  <= TRANSPORT a_N91_aIN  ;
xor2_4752: a_N91_aIN <=  n_5242  XOR n_5246;
or1_4753: n_5242 <=  n_5243;
and2_4754: n_5243 <=  n_5244  AND n_5245;
delay_4755: n_5244  <= TRANSPORT a_N1146_aOUT  ;
delay_4756: n_5245  <= TRANSPORT a_N1164_aOUT  ;
and1_4757: n_5246 <=  gnd;
delay_4758: a_LC8_D21_aOUT  <= TRANSPORT a_LC8_D21_aIN  ;
xor2_4759: a_LC8_D21_aIN <=  n_5249  XOR n_5254;
or2_4760: n_5249 <=  n_5250  OR n_5252;
and1_4761: n_5250 <=  n_5251;
delay_4762: n_5251  <= TRANSPORT a_N86_aOUT  ;
and1_4763: n_5252 <=  n_5253;
delay_4764: n_5253  <= TRANSPORT a_N91_aOUT  ;
and1_4765: n_5254 <=  gnd;
delay_4766: a_LC2_D7_aOUT  <= TRANSPORT a_LC2_D7_aIN  ;
xor2_4767: a_LC2_D7_aIN <=  n_5257  XOR n_5264;
or2_4768: n_5257 <=  n_5258  OR n_5260;
and1_4769: n_5258 <=  n_5259;
delay_4770: n_5259  <= TRANSPORT a_N1080_aOUT  ;
and3_4771: n_5260 <=  n_5261  AND n_5262  AND n_5263;
inv_4772: n_5261  <= TRANSPORT NOT a_N1175_aNOT_aOUT  ;
delay_4773: n_5262  <= TRANSPORT a_N61_aQ  ;
delay_4774: n_5263  <= TRANSPORT a_N63_aQ  ;
and1_4775: n_5264 <=  gnd;
delay_4776: a_N524_aOUT  <= TRANSPORT a_N524_aIN  ;
xor2_4777: a_N524_aIN <=  n_5267  XOR n_5277;
or3_4778: n_5267 <=  n_5268  OR n_5271  OR n_5274;
and2_4779: n_5268 <=  n_5269  AND n_5270;
inv_4780: n_5269  <= TRANSPORT NOT a_N83_aOUT  ;
delay_4781: n_5270  <= TRANSPORT a_LC8_D21_aOUT  ;
and2_4782: n_5271 <=  n_5272  AND n_5273;
inv_4783: n_5272  <= TRANSPORT NOT a_N83_aOUT  ;
delay_4784: n_5273  <= TRANSPORT a_LC2_D7_aOUT  ;
and2_4785: n_5274 <=  n_5275  AND n_5276;
inv_4786: n_5275  <= TRANSPORT NOT a_N83_aOUT  ;
inv_4787: n_5276  <= TRANSPORT NOT a_N114_aOUT  ;
and1_4788: n_5277 <=  gnd;
delay_4789: a_N1124_aNOT_aOUT  <= TRANSPORT a_N1124_aNOT_aIN  ;
xor2_4790: a_N1124_aNOT_aIN <=  n_5280  XOR n_5285;
or2_4791: n_5280 <=  n_5281  OR n_5283;
and1_4792: n_5281 <=  n_5282;
delay_4793: n_5282  <= TRANSPORT a_N676_aOUT  ;
and1_4794: n_5283 <=  n_5284;
delay_4795: n_5284  <= TRANSPORT a_N524_aOUT  ;
and1_4796: n_5285 <=  gnd;
dff_4797: DFF_a8251
    PORT MAP ( D => a_N1170_aD, CLK => a_N1170_aCLK, CLRN => a_N1170_aCLRN,
          PRN => vcc, Q => a_N1170_aQ);
delay_4798: a_N1170_aCLRN  <= TRANSPORT nRESET  ;
xor2_4799: a_N1170_aD <=  n_5292  XOR n_5306;
or3_4800: n_5292 <=  n_5293  OR n_5297  OR n_5301;
and3_4801: n_5293 <=  n_5294  AND n_5295  AND n_5296;
delay_4802: n_5294  <= TRANSPORT a_N1125_aOUT  ;
delay_4803: n_5295  <= TRANSPORT a_N1170_aQ  ;
inv_4804: n_5296  <= TRANSPORT NOT a_N1171_aQ  ;
and3_4805: n_5297 <=  n_5298  AND n_5299  AND n_5300;
delay_4806: n_5298  <= TRANSPORT a_N1125_aOUT  ;
inv_4807: n_5299  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_4808: n_5300  <= TRANSPORT a_N1170_aQ  ;
and4_4809: n_5301 <=  n_5302  AND n_5303  AND n_5304  AND n_5305;
delay_4810: n_5302  <= TRANSPORT a_N1125_aOUT  ;
delay_4811: n_5303  <= TRANSPORT a_N1124_aNOT_aOUT  ;
inv_4812: n_5304  <= TRANSPORT NOT a_N1170_aQ  ;
delay_4813: n_5305  <= TRANSPORT a_N1171_aQ  ;
and1_4814: n_5306 <=  gnd;
delay_4815: n_5307  <= TRANSPORT nRXC  ;
filter_4816: FILTER_a8251
    PORT MAP (IN1 => n_5307, Y => a_N1170_aCLK);
delay_4817: a_N376_aOUT  <= TRANSPORT a_N376_aIN  ;
xor2_4818: a_N376_aIN <=  n_5311  XOR n_5316;
or1_4819: n_5311 <=  n_5312;
and3_4820: n_5312 <=  n_5313  AND n_5314  AND n_5315;
delay_4821: n_5313  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_4822: n_5314  <= TRANSPORT a_N1170_aQ  ;
delay_4823: n_5315  <= TRANSPORT a_N1171_aQ  ;
and1_4824: n_5316 <=  gnd;
dff_4825: DFF_a8251
    PORT MAP ( D => a_N1169_aD, CLK => a_N1169_aCLK, CLRN => a_N1169_aCLRN,
          PRN => vcc, Q => a_N1169_aQ);
delay_4826: a_N1169_aCLRN  <= TRANSPORT nRESET  ;
xor2_4827: a_N1169_aD <=  n_5323  XOR n_5332;
or2_4828: n_5323 <=  n_5324  OR n_5328;
and3_4829: n_5324 <=  n_5325  AND n_5326  AND n_5327;
delay_4830: n_5325  <= TRANSPORT a_N1125_aOUT  ;
inv_4831: n_5326  <= TRANSPORT NOT a_N376_aOUT  ;
delay_4832: n_5327  <= TRANSPORT a_N1169_aQ  ;
and3_4833: n_5328 <=  n_5329  AND n_5330  AND n_5331;
delay_4834: n_5329  <= TRANSPORT a_N1125_aOUT  ;
delay_4835: n_5330  <= TRANSPORT a_N376_aOUT  ;
inv_4836: n_5331  <= TRANSPORT NOT a_N1169_aQ  ;
and1_4837: n_5332 <=  gnd;
delay_4838: n_5333  <= TRANSPORT nRXC  ;
filter_4839: FILTER_a8251
    PORT MAP (IN1 => n_5333, Y => a_N1169_aCLK);
dff_4840: DFF_a8251
    PORT MAP ( D => a_N1167_aD, CLK => a_N1167_aCLK, CLRN => a_N1167_aCLRN,
          PRN => vcc, Q => a_N1167_aQ);
delay_4841: a_N1167_aCLRN  <= TRANSPORT nRESET  ;
xor2_4842: a_N1167_aD <=  n_5341  XOR n_5355;
or3_4843: n_5341 <=  n_5342  OR n_5346  OR n_5350;
and3_4844: n_5342 <=  n_5343  AND n_5344  AND n_5345;
delay_4845: n_5343  <= TRANSPORT a_N1125_aOUT  ;
inv_4846: n_5344  <= TRANSPORT NOT a_N1169_aQ  ;
delay_4847: n_5345  <= TRANSPORT a_N1167_aQ  ;
and3_4848: n_5346 <=  n_5347  AND n_5348  AND n_5349;
delay_4849: n_5347  <= TRANSPORT a_N1125_aOUT  ;
inv_4850: n_5348  <= TRANSPORT NOT a_N376_aOUT  ;
delay_4851: n_5349  <= TRANSPORT a_N1167_aQ  ;
and4_4852: n_5350 <=  n_5351  AND n_5352  AND n_5353  AND n_5354;
delay_4853: n_5351  <= TRANSPORT a_N1125_aOUT  ;
delay_4854: n_5352  <= TRANSPORT a_N376_aOUT  ;
delay_4855: n_5353  <= TRANSPORT a_N1169_aQ  ;
inv_4856: n_5354  <= TRANSPORT NOT a_N1167_aQ  ;
and1_4857: n_5355 <=  gnd;
delay_4858: n_5356  <= TRANSPORT nRXC  ;
filter_4859: FILTER_a8251
    PORT MAP (IN1 => n_5356, Y => a_N1167_aCLK);
delay_4860: a_N720_aOUT  <= TRANSPORT a_N720_aIN  ;
xor2_4861: a_N720_aIN <=  n_5360  XOR n_5366;
or1_4862: n_5360 <=  n_5361;
and4_4863: n_5361 <=  n_5362  AND n_5363  AND n_5364  AND n_5365;
delay_4864: n_5362  <= TRANSPORT a_N1189_aOUT  ;
delay_4865: n_5363  <= TRANSPORT a_N1757_aQ  ;
delay_4866: n_5364  <= TRANSPORT a_N1756_aQ  ;
delay_4867: n_5365  <= TRANSPORT DIN(0)  ;
and1_4868: n_5366 <=  gnd;
dff_4869: DFF_a8251
    PORT MAP ( D => a_SSYNC2_F0_G_aD, CLK => a_SSYNC2_F0_G_aCLK, CLRN => a_SSYNC2_F0_G_aCLRN,
          PRN => vcc, Q => a_SSYNC2_F0_G_aQ);
delay_4870: a_SSYNC2_F0_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_4871: a_SSYNC2_F0_G_aD <=  n_5373  XOR n_5381;
or2_4872: n_5373 <=  n_5374  OR n_5378;
and3_4873: n_5374 <=  n_5375  AND n_5376  AND n_5377;
delay_4874: n_5375  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_4875: n_5376  <= TRANSPORT a_N1116_aNOT_aOUT  ;
delay_4876: n_5377  <= TRANSPORT a_SSYNC2_F0_G_aQ  ;
and2_4877: n_5378 <=  n_5379  AND n_5380;
delay_4878: n_5379  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_4879: n_5380  <= TRANSPORT a_N720_aOUT  ;
and1_4880: n_5381 <=  gnd;
delay_4881: n_5382  <= TRANSPORT CLK  ;
filter_4882: FILTER_a8251
    PORT MAP (IN1 => n_5382, Y => a_SSYNC2_F0_G_aCLK);
dff_4883: DFF_a8251
    PORT MAP ( D => a_N729_aD, CLK => a_N729_aCLK, CLRN => a_N729_aCLRN, PRN => vcc,
          Q => a_N729_aQ);
delay_4884: a_N729_aCLRN  <= TRANSPORT nRESET  ;
xor2_4885: a_N729_aD <=  n_5390  XOR n_5401;
or2_4886: n_5390 <=  n_5391  OR n_5396;
and4_4887: n_5391 <=  n_5392  AND n_5393  AND n_5394  AND n_5395;
delay_4888: n_5392  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_4889: n_5393  <= TRANSPORT a_N1032_aNOT_aOUT  ;
delay_4890: n_5394  <= TRANSPORT a_N729_aQ  ;
inv_4891: n_5395  <= TRANSPORT NOT a_SMODE_OUT_F7_G_aQ  ;
and4_4892: n_5396 <=  n_5397  AND n_5398  AND n_5399  AND n_5400;
inv_4893: n_5397  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_4894: n_5398  <= TRANSPORT a_N1032_aNOT_aOUT  ;
inv_4895: n_5399  <= TRANSPORT NOT a_N729_aQ  ;
inv_4896: n_5400  <= TRANSPORT NOT a_SMODE_OUT_F7_G_aQ  ;
and1_4897: n_5401 <=  gnd;
inv_4898: n_5402  <= TRANSPORT NOT nTXC  ;
filter_4899: FILTER_a8251
    PORT MAP (IN1 => n_5402, Y => a_N729_aCLK);
delay_4900: a_N119_aOUT  <= TRANSPORT a_N119_aIN  ;
xor2_4901: a_N119_aIN <=  n_5406  XOR n_5410;
or1_4902: n_5406 <=  n_5407;
and2_4903: n_5407 <=  n_5408  AND n_5409;
delay_4904: n_5408  <= TRANSPORT a_N1189_aOUT  ;
delay_4905: n_5409  <= TRANSPORT DIN(0)  ;
and1_4906: n_5410 <=  gnd;
dff_4907: DFF_a8251
    PORT MAP ( D => a_SSYNC1_F0_G_aD, CLK => a_SSYNC1_F0_G_aCLK, CLRN => a_SSYNC1_F0_G_aCLRN,
          PRN => vcc, Q => a_SSYNC1_F0_G_aQ);
delay_4908: a_SSYNC1_F0_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_4909: a_SSYNC1_F0_G_aD <=  n_5417  XOR n_5424;
or2_4910: n_5417 <=  n_5418  OR n_5421;
and2_4911: n_5418 <=  n_5419  AND n_5420;
delay_4912: n_5419  <= TRANSPORT a_N608_aOUT  ;
delay_4913: n_5420  <= TRANSPORT a_SSYNC1_F0_G_aQ  ;
and2_4914: n_5421 <=  n_5422  AND n_5423;
delay_4915: n_5422  <= TRANSPORT a_LC5_B5_aOUT  ;
delay_4916: n_5423  <= TRANSPORT a_N119_aOUT  ;
and1_4917: n_5424 <=  gnd;
delay_4918: n_5425  <= TRANSPORT CLK  ;
filter_4919: FILTER_a8251
    PORT MAP (IN1 => n_5425, Y => a_SSYNC1_F0_G_aCLK);
dff_4920: DFF_a8251
    PORT MAP ( D => a_N2030_aD, CLK => a_N2030_aCLK, CLRN => a_N2030_aCLRN,
          PRN => vcc, Q => a_N2030_aQ);
delay_4921: a_N2030_aCLRN  <= TRANSPORT nRESET  ;
xor2_4922: a_N2030_aD <=  n_5434  XOR n_5441;
or2_4923: n_5434 <=  n_5435  OR n_5438;
and2_4924: n_5435 <=  n_5436  AND n_5437;
delay_4925: n_5436  <= TRANSPORT a_N1198_aOUT  ;
delay_4926: n_5437  <= TRANSPORT a_N2030_aQ  ;
and2_4927: n_5438 <=  n_5439  AND n_5440;
delay_4928: n_5439  <= TRANSPORT a_N1197_aOUT  ;
delay_4929: n_5440  <= TRANSPORT DIN(1)  ;
and1_4930: n_5441 <=  gnd;
inv_4931: n_5442  <= TRANSPORT NOT nTXC  ;
filter_4932: FILTER_a8251
    PORT MAP (IN1 => n_5442, Y => a_N2030_aCLK);
dff_4933: DFF_a8251
    PORT MAP ( D => a_N2029_aD, CLK => a_N2029_aCLK, CLRN => a_N2029_aCLRN,
          PRN => vcc, Q => a_N2029_aQ);
delay_4934: a_N2029_aCLRN  <= TRANSPORT nRESET  ;
xor2_4935: a_N2029_aD <=  n_5450  XOR n_5457;
or2_4936: n_5450 <=  n_5451  OR n_5454;
and2_4937: n_5451 <=  n_5452  AND n_5453;
delay_4938: n_5452  <= TRANSPORT a_N1197_aOUT  ;
delay_4939: n_5453  <= TRANSPORT DIN(2)  ;
and2_4940: n_5454 <=  n_5455  AND n_5456;
delay_4941: n_5455  <= TRANSPORT a_N1198_aOUT  ;
delay_4942: n_5456  <= TRANSPORT a_N2029_aQ  ;
and1_4943: n_5457 <=  gnd;
inv_4944: n_5458  <= TRANSPORT NOT nTXC  ;
filter_4945: FILTER_a8251
    PORT MAP (IN1 => n_5458, Y => a_N2029_aCLK);
dff_4946: DFF_a8251
    PORT MAP ( D => a_N2028_aD, CLK => a_N2028_aCLK, CLRN => a_N2028_aCLRN,
          PRN => vcc, Q => a_N2028_aQ);
delay_4947: a_N2028_aCLRN  <= TRANSPORT nRESET  ;
xor2_4948: a_N2028_aD <=  n_5466  XOR n_5473;
or2_4949: n_5466 <=  n_5467  OR n_5470;
and2_4950: n_5467 <=  n_5468  AND n_5469;
delay_4951: n_5468  <= TRANSPORT a_N1198_aOUT  ;
delay_4952: n_5469  <= TRANSPORT a_N2028_aQ  ;
and2_4953: n_5470 <=  n_5471  AND n_5472;
delay_4954: n_5471  <= TRANSPORT a_N1197_aOUT  ;
delay_4955: n_5472  <= TRANSPORT DIN(3)  ;
and1_4956: n_5473 <=  gnd;
inv_4957: n_5474  <= TRANSPORT NOT nTXC  ;
filter_4958: FILTER_a8251
    PORT MAP (IN1 => n_5474, Y => a_N2028_aCLK);
delay_4959: a_LC2_B1_aOUT  <= TRANSPORT a_LC2_B1_aIN  ;
xor2_4960: a_LC2_B1_aIN <=  n_5478  XOR n_5484;
or1_4961: n_5478 <=  n_5479;
and4_4962: n_5479 <=  n_5480  AND n_5481  AND n_5482  AND n_5483;
inv_4963: n_5480  <= TRANSPORT NOT a_LC7_B6_aNOT_aOUT  ;
delay_4964: n_5481  <= TRANSPORT a_N362_aQ  ;
delay_4965: n_5482  <= TRANSPORT a_N360_aQ  ;
delay_4966: n_5483  <= TRANSPORT a_N361_aQ  ;
and1_4967: n_5484 <=  gnd;
dff_4968: DFF_a8251
    PORT MAP ( D => a_N359_aD, CLK => a_N359_aCLK, CLRN => a_N359_aCLRN, PRN => vcc,
          Q => a_N359_aQ);
delay_4969: a_N359_aCLRN  <= TRANSPORT nRESET  ;
xor2_4970: a_N359_aD <=  n_5491  XOR n_5503;
or3_4971: n_5491 <=  n_5492  OR n_5496  OR n_5500;
and3_4972: n_5492 <=  n_5493  AND n_5494  AND n_5495;
delay_4973: n_5493  <= TRANSPORT a_LC4_B10_aOUT  ;
inv_4974: n_5494  <= TRANSPORT NOT a_LC2_B1_aOUT  ;
delay_4975: n_5495  <= TRANSPORT a_N359_aQ  ;
and3_4976: n_5496 <=  n_5497  AND n_5498  AND n_5499;
delay_4977: n_5497  <= TRANSPORT a_LC4_B10_aOUT  ;
delay_4978: n_5498  <= TRANSPORT a_LC2_B1_aOUT  ;
inv_4979: n_5499  <= TRANSPORT NOT a_N359_aQ  ;
and2_4980: n_5500 <=  n_5501  AND n_5502;
delay_4981: n_5501  <= TRANSPORT a_LC1_B10_aOUT  ;
delay_4982: n_5502  <= TRANSPORT a_N359_aQ  ;
and1_4983: n_5503 <=  gnd;
inv_4984: n_5504  <= TRANSPORT NOT nTXC  ;
filter_4985: FILTER_a8251
    PORT MAP (IN1 => n_5504, Y => a_N359_aCLK);
dff_4986: DFF_a8251
    PORT MAP ( D => a_N396_aD, CLK => a_N396_aCLK, CLRN => a_N396_aCLRN, PRN => vcc,
          Q => a_N396_aQ);
delay_4987: a_N396_aCLRN  <= TRANSPORT nRESET  ;
xor2_4988: a_N396_aD <=  n_5512  XOR n_5526;
or3_4989: n_5512 <=  n_5513  OR n_5517  OR n_5521;
and3_4990: n_5513 <=  n_5514  AND n_5515  AND n_5516;
delay_4991: n_5514  <= TRANSPORT a_N1056_aOUT  ;
delay_4992: n_5515  <= TRANSPORT a_N396_aQ  ;
inv_4993: n_5516  <= TRANSPORT NOT a_N397_aQ  ;
and3_4994: n_5517 <=  n_5518  AND n_5519  AND n_5520;
delay_4995: n_5518  <= TRANSPORT a_N470_aOUT  ;
delay_4996: n_5519  <= TRANSPORT a_N1056_aOUT  ;
delay_4997: n_5520  <= TRANSPORT a_N396_aQ  ;
and4_4998: n_5521 <=  n_5522  AND n_5523  AND n_5524  AND n_5525;
inv_4999: n_5522  <= TRANSPORT NOT a_N470_aOUT  ;
delay_5000: n_5523  <= TRANSPORT a_N1056_aOUT  ;
inv_5001: n_5524  <= TRANSPORT NOT a_N396_aQ  ;
delay_5002: n_5525  <= TRANSPORT a_N397_aQ  ;
and1_5003: n_5526 <=  gnd;
inv_5004: n_5527  <= TRANSPORT NOT nTXC  ;
filter_5005: FILTER_a8251
    PORT MAP (IN1 => n_5527, Y => a_N396_aCLK);
dff_5006: DFF_a8251
    PORT MAP ( D => a_N397_aD, CLK => a_N397_aCLK, CLRN => a_N397_aCLRN, PRN => vcc,
          Q => a_N397_aQ);
delay_5007: a_N397_aCLRN  <= TRANSPORT nRESET  ;
xor2_5008: a_N397_aD <=  n_5535  XOR n_5544;
or2_5009: n_5535 <=  n_5536  OR n_5540;
and3_5010: n_5536 <=  n_5537  AND n_5538  AND n_5539;
inv_5011: n_5537  <= TRANSPORT NOT a_N470_aOUT  ;
delay_5012: n_5538  <= TRANSPORT a_N1056_aOUT  ;
inv_5013: n_5539  <= TRANSPORT NOT a_N397_aQ  ;
and3_5014: n_5540 <=  n_5541  AND n_5542  AND n_5543;
delay_5015: n_5541  <= TRANSPORT a_N470_aOUT  ;
delay_5016: n_5542  <= TRANSPORT a_N1056_aOUT  ;
delay_5017: n_5543  <= TRANSPORT a_N397_aQ  ;
and1_5018: n_5544 <=  gnd;
inv_5019: n_5545  <= TRANSPORT NOT nTXC  ;
filter_5020: FILTER_a8251
    PORT MAP (IN1 => n_5545, Y => a_N397_aCLK);
dff_5021: DFF_a8251
    PORT MAP ( D => a_N1171_aD, CLK => a_N1171_aCLK, CLRN => a_N1171_aCLRN,
          PRN => vcc, Q => a_N1171_aQ);
delay_5022: a_N1171_aCLRN  <= TRANSPORT nRESET  ;
xor2_5023: a_N1171_aD <=  n_5553  XOR n_5562;
or2_5024: n_5553 <=  n_5554  OR n_5558;
and3_5025: n_5554 <=  n_5555  AND n_5556  AND n_5557;
delay_5026: n_5555  <= TRANSPORT a_N1125_aOUT  ;
inv_5027: n_5556  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5028: n_5557  <= TRANSPORT a_N1171_aQ  ;
and3_5029: n_5558 <=  n_5559  AND n_5560  AND n_5561;
delay_5030: n_5559  <= TRANSPORT a_N1125_aOUT  ;
delay_5031: n_5560  <= TRANSPORT a_N1124_aNOT_aOUT  ;
inv_5032: n_5561  <= TRANSPORT NOT a_N1171_aQ  ;
and1_5033: n_5562 <=  gnd;
delay_5034: n_5563  <= TRANSPORT nRXC  ;
filter_5035: FILTER_a8251
    PORT MAP (IN1 => n_5563, Y => a_N1171_aCLK);
delay_5036: a_LC3_A3_aOUT  <= TRANSPORT a_LC3_A3_aIN  ;
xor2_5037: a_LC3_A3_aIN <=  n_5567  XOR n_5573;
or1_5038: n_5567 <=  n_5568;
and3_5039: n_5568 <=  n_5569  AND n_5571  AND n_5572;
delay_5040: n_5569  <= TRANSPORT a_N1553_aQ  ;
inv_5041: n_5571  <= TRANSPORT NOT a_N1555_aQ  ;
inv_5042: n_5572  <= TRANSPORT NOT a_N1556_aQ  ;
and1_5043: n_5573 <=  gnd;
delay_5044: a_LC3_D4_aNOT_aOUT  <= TRANSPORT a_LC3_D4_aNOT_aIN  ;
xor2_5045: a_LC3_D4_aNOT_aIN <=  n_5576  XOR n_5582;
or1_5046: n_5576 <=  n_5577;
and4_5047: n_5577 <=  n_5578  AND n_5579  AND n_5580  AND n_5581;
delay_5048: n_5578  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5049: n_5579  <= TRANSPORT a_N64_aQ  ;
inv_5050: n_5580  <= TRANSPORT NOT a_N61_aQ  ;
inv_5051: n_5581  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and1_5052: n_5582 <=  gnd;
delay_5053: a_LC4_D4_aOUT  <= TRANSPORT a_LC4_D4_aIN  ;
xor2_5054: a_LC4_D4_aIN <=  n_5585  XOR n_5590;
or1_5055: n_5585 <=  n_5586;
and3_5056: n_5586 <=  n_5587  AND n_5588  AND n_5589;
inv_5057: n_5587  <= TRANSPORT NOT a_N132_aOUT  ;
delay_5058: n_5588  <= TRANSPORT a_N1146_aOUT  ;
delay_5059: n_5589  <= TRANSPORT a_LC3_D4_aNOT_aOUT  ;
and1_5060: n_5590 <=  gnd;
delay_5061: a_LC2_D4_aOUT  <= TRANSPORT a_LC2_D4_aIN  ;
xor2_5062: a_LC2_D4_aIN <=  n_5593  XOR n_5599;
or1_5063: n_5593 <=  n_5594;
and4_5064: n_5594 <=  n_5595  AND n_5596  AND n_5597  AND n_5598;
delay_5065: n_5595  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5066: n_5596  <= TRANSPORT a_N127_aOUT  ;
delay_5067: n_5597  <= TRANSPORT a_N62_aQ  ;
inv_5068: n_5598  <= TRANSPORT NOT a_N63_aQ  ;
and1_5069: n_5599 <=  gnd;
delay_5070: a_LC5_D4_aOUT  <= TRANSPORT a_LC5_D4_aIN  ;
xor2_5071: a_LC5_D4_aIN <=  n_5602  XOR n_5608;
or1_5072: n_5602 <=  n_5603;
and4_5073: n_5603 <=  n_5604  AND n_5605  AND n_5606  AND n_5607;
delay_5074: n_5604  <= TRANSPORT a_N1183_aNOT_aOUT  ;
delay_5075: n_5605  <= TRANSPORT a_N1164_aOUT  ;
delay_5076: n_5606  <= TRANSPORT a_N62_aQ  ;
inv_5077: n_5607  <= TRANSPORT NOT a_N63_aQ  ;
and1_5078: n_5608 <=  gnd;
delay_5079: a_LC6_D4_aOUT  <= TRANSPORT a_LC6_D4_aIN  ;
xor2_5080: a_LC6_D4_aIN <=  n_5610  XOR n_5619;
or3_5081: n_5610 <=  n_5611  OR n_5614  OR n_5617;
and2_5082: n_5611 <=  n_5612  AND n_5613;
delay_5083: n_5612  <= TRANSPORT a_LC4_D4_aOUT  ;
delay_5084: n_5613  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and2_5085: n_5614 <=  n_5615  AND n_5616;
delay_5086: n_5615  <= TRANSPORT a_LC2_D4_aOUT  ;
delay_5087: n_5616  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_5088: n_5617 <=  n_5618;
delay_5089: n_5618  <= TRANSPORT a_LC5_D4_aOUT  ;
and1_5090: n_5619 <=  gnd;
delay_5091: a_N1145_aOUT  <= TRANSPORT a_N1145_aIN  ;
xor2_5092: a_N1145_aIN <=  n_5621  XOR n_5626;
or1_5093: n_5621 <=  n_5622;
and3_5094: n_5622 <=  n_5623  AND n_5624  AND n_5625;
delay_5095: n_5623  <= TRANSPORT a_N59_aQ  ;
inv_5096: n_5624  <= TRANSPORT NOT a_N62_aQ  ;
inv_5097: n_5625  <= TRANSPORT NOT a_N61_aQ  ;
and1_5098: n_5626 <=  gnd;
delay_5099: a_N467_aNOT_aOUT  <= TRANSPORT a_N467_aNOT_aIN  ;
xor2_5100: a_N467_aNOT_aIN <=  n_5629  XOR n_5639;
or2_5101: n_5629 <=  n_5630  OR n_5634;
and3_5102: n_5630 <=  n_5631  AND n_5632  AND n_5633;
delay_5103: n_5631  <= TRANSPORT a_N1145_aOUT  ;
inv_5104: n_5632  <= TRANSPORT NOT a_N64_aQ  ;
delay_5105: n_5633  <= TRANSPORT a_N63_aQ  ;
and4_5106: n_5634 <=  n_5635  AND n_5636  AND n_5637  AND n_5638;
delay_5107: n_5635  <= TRANSPORT a_N1183_aNOT_aOUT  ;
delay_5108: n_5636  <= TRANSPORT a_N1145_aOUT  ;
delay_5109: n_5637  <= TRANSPORT a_N64_aQ  ;
inv_5110: n_5638  <= TRANSPORT NOT a_N63_aQ  ;
and1_5111: n_5639 <=  gnd;
delay_5112: a_N113_aNOT_aOUT  <= TRANSPORT a_N113_aNOT_aIN  ;
xor2_5113: a_N113_aNOT_aIN <=  n_5642  XOR n_5649;
or2_5114: n_5642 <=  n_5643  OR n_5645;
and1_5115: n_5643 <=  n_5644;
delay_5116: n_5644  <= TRANSPORT a_N467_aNOT_aOUT  ;
and3_5117: n_5645 <=  n_5646  AND n_5647  AND n_5648;
inv_5118: n_5646  <= TRANSPORT NOT a_N1137_aNOT_aOUT  ;
delay_5119: n_5647  <= TRANSPORT a_N61_aQ  ;
delay_5120: n_5648  <= TRANSPORT a_N63_aQ  ;
and1_5121: n_5649 <=  gnd;
delay_5122: a_N79_aNOT_aOUT  <= TRANSPORT a_N79_aNOT_aIN  ;
xor2_5123: a_N79_aNOT_aIN <=  n_5651  XOR n_5656;
or2_5124: n_5651 <=  n_5652  OR n_5654;
and1_5125: n_5652 <=  n_5653;
delay_5126: n_5653  <= TRANSPORT a_LC6_D4_aOUT  ;
and1_5127: n_5654 <=  n_5655;
delay_5128: n_5655  <= TRANSPORT a_N113_aNOT_aOUT  ;
and1_5129: n_5656 <=  gnd;
delay_5130: a_LC2_A3_aOUT  <= TRANSPORT a_LC2_A3_aIN  ;
xor2_5131: a_LC2_A3_aIN <=  n_5659  XOR n_5666;
or2_5132: n_5659 <=  n_5660  OR n_5663;
and2_5133: n_5660 <=  n_5661  AND n_5662;
delay_5134: n_5661  <= TRANSPORT a_LC3_A3_aOUT  ;
inv_5135: n_5662  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
and2_5136: n_5663 <=  n_5664  AND n_5665;
delay_5137: n_5664  <= TRANSPORT a_N1194_aNOT_aOUT  ;
delay_5138: n_5665  <= TRANSPORT a_LC3_A3_aOUT  ;
and1_5139: n_5666 <=  gnd;
delay_5140: a_N1160_aOUT  <= TRANSPORT a_N1160_aIN  ;
xor2_5141: a_N1160_aIN <=  n_5669  XOR n_5673;
or1_5142: n_5669 <=  n_5670;
and2_5143: n_5670 <=  n_5671  AND n_5672;
delay_5144: n_5671  <= TRANSPORT a_N1555_aQ  ;
delay_5145: n_5672  <= TRANSPORT a_N1556_aQ  ;
and1_5146: n_5673 <=  gnd;
delay_5147: a_N1117_aOUT  <= TRANSPORT a_N1117_aIN  ;
xor2_5148: a_N1117_aIN <=  n_5676  XOR n_5680;
or1_5149: n_5676 <=  n_5677;
and2_5150: n_5677 <=  n_5678  AND n_5679;
inv_5151: n_5678  <= TRANSPORT NOT a_N135_aOUT  ;
inv_5152: n_5679  <= TRANSPORT NOT a_SMODE_OUT_F7_G_aQ  ;
and1_5153: n_5680 <=  gnd;
delay_5154: a_LC6_A3_aOUT  <= TRANSPORT a_LC6_A3_aIN  ;
xor2_5155: a_LC6_A3_aIN <=  n_5683  XOR n_5688;
or1_5156: n_5683 <=  n_5684;
and3_5157: n_5684 <=  n_5685  AND n_5686  AND n_5687;
delay_5158: n_5685  <= TRANSPORT a_N79_aNOT_aOUT  ;
delay_5159: n_5686  <= TRANSPORT a_N1160_aOUT  ;
delay_5160: n_5687  <= TRANSPORT a_N1117_aOUT  ;
and1_5161: n_5688 <=  gnd;
dff_5162: DFF_a8251
    PORT MAP ( D => a_N1553_aD, CLK => a_N1553_aCLK, CLRN => a_N1553_aCLRN,
          PRN => vcc, Q => a_N1553_aQ);
delay_5163: a_N1553_aCLRN  <= TRANSPORT nRESET  ;
xor2_5164: a_N1553_aD <=  n_5695  XOR n_5704;
or2_5165: n_5695 <=  n_5696  OR n_5700;
and3_5166: n_5696 <=  n_5697  AND n_5698  AND n_5699;
delay_5167: n_5697  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5168: n_5698  <= TRANSPORT a_N1187_aOUT  ;
delay_5169: n_5699  <= TRANSPORT a_LC2_A3_aOUT  ;
and3_5170: n_5700 <=  n_5701  AND n_5702  AND n_5703;
delay_5171: n_5701  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5172: n_5702  <= TRANSPORT a_N1187_aOUT  ;
delay_5173: n_5703  <= TRANSPORT a_LC6_A3_aOUT  ;
and1_5174: n_5704 <=  gnd;
delay_5175: n_5705  <= TRANSPORT nRXC  ;
filter_5176: FILTER_a8251
    PORT MAP (IN1 => n_5705, Y => a_N1553_aCLK);
dff_5177: DFF_a8251
    PORT MAP ( D => a_N1307_aD, CLK => a_N1307_aCLK, CLRN => a_N1307_aCLRN,
          PRN => vcc, Q => a_N1307_aQ);
delay_5178: a_N1307_aCLRN  <= TRANSPORT nRESET  ;
xor2_5179: a_N1307_aD <=  n_5713  XOR n_5722;
or2_5180: n_5713 <=  n_5714  OR n_5718;
and3_5181: n_5714 <=  n_5715  AND n_5716  AND n_5717;
inv_5182: n_5715  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5183: n_5716  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5184: n_5717  <= TRANSPORT a_N1307_aQ  ;
and3_5185: n_5718 <=  n_5719  AND n_5720  AND n_5721;
inv_5186: n_5719  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5187: n_5720  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5188: n_5721  <= TRANSPORT a_N1306_aQ  ;
and1_5189: n_5722 <=  gnd;
delay_5190: n_5723  <= TRANSPORT nRXC  ;
filter_5191: FILTER_a8251
    PORT MAP (IN1 => n_5723, Y => a_N1307_aCLK);
dff_5192: DFF_a8251
    PORT MAP ( D => a_N1306_aD, CLK => a_N1306_aCLK, CLRN => a_N1306_aCLRN,
          PRN => vcc, Q => a_N1306_aQ);
delay_5193: a_N1306_aCLRN  <= TRANSPORT nRESET  ;
xor2_5194: a_N1306_aD <=  n_5731  XOR n_5740;
or2_5195: n_5731 <=  n_5732  OR n_5736;
and3_5196: n_5732 <=  n_5733  AND n_5734  AND n_5735;
inv_5197: n_5733  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5198: n_5734  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5199: n_5735  <= TRANSPORT a_N1306_aQ  ;
and3_5200: n_5736 <=  n_5737  AND n_5738  AND n_5739;
inv_5201: n_5737  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5202: n_5738  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5203: n_5739  <= TRANSPORT a_N1305_aQ  ;
and1_5204: n_5740 <=  gnd;
delay_5205: n_5741  <= TRANSPORT nRXC  ;
filter_5206: FILTER_a8251
    PORT MAP (IN1 => n_5741, Y => a_N1306_aCLK);
delay_5207: a_N1069_aOUT  <= TRANSPORT a_N1069_aIN  ;
xor2_5208: a_N1069_aIN <=  n_5745  XOR n_5751;
or1_5209: n_5745 <=  n_5746;
and4_5210: n_5746 <=  n_5747  AND n_5748  AND n_5749  AND n_5750;
inv_5211: n_5747  <= TRANSPORT NOT a_N1183_aNOT_aOUT  ;
delay_5212: n_5748  <= TRANSPORT a_N1145_aOUT  ;
delay_5213: n_5749  <= TRANSPORT a_N64_aQ  ;
inv_5214: n_5750  <= TRANSPORT NOT a_N63_aQ  ;
and1_5215: n_5751 <=  gnd;
dff_5216: DFF_a8251
    PORT MAP ( D => a_N59_aD, CLK => a_N59_aCLK, CLRN => a_N59_aCLRN, PRN => vcc,
          Q => a_N59_aQ);
delay_5217: a_N59_aCLRN  <= TRANSPORT nRESET  ;
xor2_5218: a_N59_aD <=  n_5758  XOR n_5768;
or3_5219: n_5758 <=  n_5759  OR n_5762  OR n_5765;
and2_5220: n_5759 <=  n_5760  AND n_5761;
inv_5221: n_5760  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5222: n_5761  <= TRANSPORT a_N1069_aOUT  ;
and2_5223: n_5762 <=  n_5763  AND n_5764;
inv_5224: n_5763  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5225: n_5764  <= TRANSPORT a_N86_aOUT  ;
and2_5226: n_5765 <=  n_5766  AND n_5767;
inv_5227: n_5766  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5228: n_5767  <= TRANSPORT NOT a_N1072_aNOT_aOUT  ;
and1_5229: n_5768 <=  gnd;
delay_5230: n_5769  <= TRANSPORT nRXC  ;
filter_5231: FILTER_a8251
    PORT MAP (IN1 => n_5769, Y => a_N59_aCLK);
dff_5232: DFF_a8251
    PORT MAP ( D => a_N1302_aD, CLK => a_N1302_aCLK, CLRN => a_N1302_aCLRN,
          PRN => vcc, Q => a_N1302_aQ);
delay_5233: a_N1302_aCLRN  <= TRANSPORT nRESET  ;
xor2_5234: a_N1302_aD <=  n_5777  XOR n_5786;
or2_5235: n_5777 <=  n_5778  OR n_5782;
and3_5236: n_5778 <=  n_5779  AND n_5780  AND n_5781;
inv_5237: n_5779  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5238: n_5780  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5239: n_5781  <= TRANSPORT a_N1301_aQ  ;
and3_5240: n_5782 <=  n_5783  AND n_5784  AND n_5785;
inv_5241: n_5783  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5242: n_5784  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5243: n_5785  <= TRANSPORT a_N1302_aQ  ;
and1_5244: n_5786 <=  gnd;
delay_5245: n_5787  <= TRANSPORT nRXC  ;
filter_5246: FILTER_a8251
    PORT MAP (IN1 => n_5787, Y => a_N1302_aCLK);
delay_5247: a_LC4_B18_aOUT  <= TRANSPORT a_LC4_B18_aIN  ;
xor2_5248: a_LC4_B18_aIN <=  n_5791  XOR n_5798;
or2_5249: n_5791 <=  n_5792  OR n_5795;
and2_5250: n_5792 <=  n_5793  AND n_5794;
delay_5251: n_5793  <= TRANSPORT a_N470_aOUT  ;
delay_5252: n_5794  <= TRANSPORT a_N606_aQ  ;
and2_5253: n_5795 <=  n_5796  AND n_5797;
delay_5254: n_5796  <= TRANSPORT a_LC2_B11_aOUT  ;
delay_5255: n_5797  <= TRANSPORT a_N605_aQ  ;
and1_5256: n_5798 <=  gnd;
delay_5257: a_N178_aOUT  <= TRANSPORT a_N178_aIN  ;
xor2_5258: a_N178_aIN <=  n_5801  XOR n_5808;
or2_5259: n_5801 <=  n_5802  OR n_5805;
and2_5260: n_5802 <=  n_5803  AND n_5804;
delay_5261: n_5803  <= TRANSPORT a_SSYNC1_F1_G_aQ  ;
inv_5262: n_5804  <= TRANSPORT NOT a_N729_aQ  ;
and2_5263: n_5805 <=  n_5806  AND n_5807;
delay_5264: n_5806  <= TRANSPORT a_SSYNC2_F1_G_aQ  ;
delay_5265: n_5807  <= TRANSPORT a_N729_aQ  ;
and1_5266: n_5808 <=  gnd;
delay_5267: a_N1094_aNOT_aOUT  <= TRANSPORT a_N1094_aNOT_aIN  ;
xor2_5268: a_N1094_aNOT_aIN <=  n_5810  XOR n_5817;
or2_5269: n_5810 <=  n_5811  OR n_5814;
and2_5270: n_5811 <=  n_5812  AND n_5813;
inv_5271: n_5812  <= TRANSPORT NOT a_N1114_aNOT_aOUT  ;
delay_5272: n_5813  <= TRANSPORT a_N178_aOUT  ;
and2_5273: n_5814 <=  n_5815  AND n_5816;
delay_5274: n_5815  <= TRANSPORT a_N1114_aNOT_aOUT  ;
delay_5275: n_5816  <= TRANSPORT a_N2030_aQ  ;
and1_5276: n_5817 <=  gnd;
dff_5277: DFF_a8251
    PORT MAP ( D => a_N606_aD, CLK => a_N606_aCLK, CLRN => a_N606_aCLRN, PRN => vcc,
          Q => a_N606_aQ);
delay_5278: a_N606_aCLRN  <= TRANSPORT nRESET  ;
xor2_5279: a_N606_aD <=  n_5824  XOR n_5833;
or2_5280: n_5824 <=  n_5825  OR n_5829;
and3_5281: n_5825 <=  n_5826  AND n_5827  AND n_5828;
delay_5282: n_5826  <= TRANSPORT a_N81_aNOT_aOUT  ;
delay_5283: n_5827  <= TRANSPORT a_N221_aNOT_aOUT  ;
delay_5284: n_5828  <= TRANSPORT a_LC4_B18_aOUT  ;
and3_5285: n_5829 <=  n_5830  AND n_5831  AND n_5832;
delay_5286: n_5830  <= TRANSPORT a_N81_aNOT_aOUT  ;
inv_5287: n_5831  <= TRANSPORT NOT a_N221_aNOT_aOUT  ;
delay_5288: n_5832  <= TRANSPORT a_N1094_aNOT_aOUT  ;
and1_5289: n_5833 <=  gnd;
inv_5290: n_5834  <= TRANSPORT NOT nTXC  ;
filter_5291: FILTER_a8251
    PORT MAP (IN1 => n_5834, Y => a_N606_aCLK);
delay_5292: a_LC4_A7_aOUT  <= TRANSPORT a_LC4_A7_aIN  ;
xor2_5293: a_LC4_A7_aIN <=  n_5838  XOR n_5848;
or2_5294: n_5838 <=  n_5839  OR n_5843;
and3_5295: n_5839 <=  n_5840  AND n_5841  AND n_5842;
delay_5296: n_5840  <= TRANSPORT a_N1117_aOUT  ;
inv_5297: n_5841  <= TRANSPORT NOT a_N1555_aQ  ;
delay_5298: n_5842  <= TRANSPORT a_N1556_aQ  ;
and4_5299: n_5843 <=  n_5844  AND n_5845  AND n_5846  AND n_5847;
delay_5300: n_5844  <= TRANSPORT a_N1120_aNOT_aOUT  ;
inv_5301: n_5845  <= TRANSPORT NOT a_N1117_aOUT  ;
delay_5302: n_5846  <= TRANSPORT a_N1555_aQ  ;
delay_5303: n_5847  <= TRANSPORT a_N1556_aQ  ;
and1_5304: n_5848 <=  gnd;
delay_5305: a_LC2_A7_aOUT  <= TRANSPORT a_LC2_A7_aIN  ;
xor2_5306: a_LC2_A7_aIN <=  n_5851  XOR n_5860;
or2_5307: n_5851 <=  n_5852  OR n_5856;
and3_5308: n_5852 <=  n_5853  AND n_5854  AND n_5855;
inv_5309: n_5853  <= TRANSPORT NOT a_N1194_aNOT_aOUT  ;
delay_5310: n_5854  <= TRANSPORT a_N1555_aQ  ;
inv_5311: n_5855  <= TRANSPORT NOT a_N1556_aQ  ;
and3_5312: n_5856 <=  n_5857  AND n_5858  AND n_5859;
delay_5313: n_5857  <= TRANSPORT a_N132_aOUT  ;
delay_5314: n_5858  <= TRANSPORT a_N1555_aQ  ;
inv_5315: n_5859  <= TRANSPORT NOT a_N1556_aQ  ;
and1_5316: n_5860 <=  gnd;
delay_5317: a_N134_aNOT_aOUT  <= TRANSPORT a_N134_aNOT_aIN  ;
xor2_5318: a_N134_aNOT_aIN <=  n_5862  XOR n_5866;
or1_5319: n_5862 <=  n_5863;
and2_5320: n_5863 <=  n_5864  AND n_5865;
inv_5321: n_5864  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5322: n_5865  <= TRANSPORT a_N79_aNOT_aOUT  ;
and1_5323: n_5866 <=  gnd;
delay_5324: a_N1193_aOUT  <= TRANSPORT a_N1193_aIN  ;
xor2_5325: a_N1193_aIN <=  n_5869  XOR n_5874;
or1_5326: n_5869 <=  n_5870;
and3_5327: n_5870 <=  n_5871  AND n_5872  AND n_5873;
inv_5328: n_5871  <= TRANSPORT NOT a_N1194_aNOT_aOUT  ;
delay_5329: n_5872  <= TRANSPORT a_LC3_A3_aOUT  ;
delay_5330: n_5873  <= TRANSPORT a_N134_aNOT_aOUT  ;
and1_5331: n_5874 <=  gnd;
delay_5332: a_N278_aOUT  <= TRANSPORT a_N278_aIN  ;
xor2_5333: a_N278_aIN <=  n_5877  XOR n_5885;
or2_5334: n_5877 <=  n_5878  OR n_5881;
and2_5335: n_5878 <=  n_5879  AND n_5880;
delay_5336: n_5879  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5337: n_5880  <= TRANSPORT a_N1193_aOUT  ;
and3_5338: n_5881 <=  n_5882  AND n_5883  AND n_5884;
delay_5339: n_5882  <= TRANSPORT a_N1120_aNOT_aOUT  ;
inv_5340: n_5883  <= TRANSPORT NOT a_N79_aNOT_aOUT  ;
delay_5341: n_5884  <= TRANSPORT a_N1160_aOUT  ;
and1_5342: n_5885 <=  gnd;
delay_5343: a_LC6_A13_aOUT  <= TRANSPORT a_LC6_A13_aIN  ;
xor2_5344: a_LC6_A13_aIN <=  n_5888  XOR n_5893;
or1_5345: n_5888 <=  n_5889;
and3_5346: n_5889 <=  n_5890  AND n_5891  AND n_5892;
inv_5347: n_5890  <= TRANSPORT NOT a_N135_aOUT  ;
delay_5348: n_5891  <= TRANSPORT a_N1556_aQ  ;
delay_5349: n_5892  <= TRANSPORT a_SMODE_OUT_F7_G_aQ  ;
and1_5350: n_5893 <=  gnd;
delay_5351: a_LC2_A13_aOUT  <= TRANSPORT a_LC2_A13_aIN  ;
xor2_5352: a_LC2_A13_aIN <=  n_5896  XOR n_5905;
or3_5353: n_5896 <=  n_5897  OR n_5900  OR n_5903;
and2_5354: n_5897 <=  n_5898  AND n_5899;
delay_5355: n_5898  <= TRANSPORT a_LC6_A13_aOUT  ;
inv_5356: n_5899  <= TRANSPORT NOT a_N1555_aQ  ;
and2_5357: n_5900 <=  n_5901  AND n_5902;
delay_5358: n_5901  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5359: n_5902  <= TRANSPORT a_LC6_A13_aOUT  ;
and1_5360: n_5903 <=  n_5904;
inv_5361: n_5904  <= TRANSPORT NOT a_N1037_aNOT_aOUT  ;
and1_5362: n_5905 <=  gnd;
delay_5363: a_N264_aNOT_aOUT  <= TRANSPORT a_N264_aNOT_aIN  ;
xor2_5364: a_N264_aNOT_aIN <=  n_5908  XOR n_5917;
or2_5365: n_5908 <=  n_5909  OR n_5913;
and3_5366: n_5909 <=  n_5910  AND n_5911  AND n_5912;
delay_5367: n_5910  <= TRANSPORT a_N1187_aOUT  ;
delay_5368: n_5911  <= TRANSPORT a_N278_aOUT  ;
delay_5369: n_5912  <= TRANSPORT nRESET  ;
and3_5370: n_5913 <=  n_5914  AND n_5915  AND n_5916;
delay_5371: n_5914  <= TRANSPORT a_N1187_aOUT  ;
delay_5372: n_5915  <= TRANSPORT a_LC2_A13_aOUT  ;
delay_5373: n_5916  <= TRANSPORT nRESET  ;
and1_5374: n_5917 <=  gnd;
dff_5375: DFF_a8251
    PORT MAP ( D => a_N1555_aD, CLK => a_N1555_aCLK, CLRN => a_N1555_aCLRN,
          PRN => vcc, Q => a_N1555_aQ);
delay_5376: a_N1555_aCLRN  <= TRANSPORT nRESET  ;
xor2_5377: a_N1555_aD <=  n_5924  XOR n_5933;
or3_5378: n_5924 <=  n_5925  OR n_5928  OR n_5931;
and2_5379: n_5925 <=  n_5926  AND n_5927;
delay_5380: n_5926  <= TRANSPORT a_N1187_aOUT  ;
delay_5381: n_5927  <= TRANSPORT a_LC4_A7_aOUT  ;
and2_5382: n_5928 <=  n_5929  AND n_5930;
delay_5383: n_5929  <= TRANSPORT a_N1187_aOUT  ;
delay_5384: n_5930  <= TRANSPORT a_LC2_A7_aOUT  ;
and1_5385: n_5931 <=  n_5932;
delay_5386: n_5932  <= TRANSPORT a_N264_aNOT_aOUT  ;
and1_5387: n_5933 <=  gnd;
delay_5388: n_5934  <= TRANSPORT nRXC  ;
filter_5389: FILTER_a8251
    PORT MAP (IN1 => n_5934, Y => a_N1555_aCLK);
delay_5390: a_LC4_A3_aOUT  <= TRANSPORT a_LC4_A3_aIN  ;
xor2_5391: a_LC4_A3_aIN <=  n_5938  XOR n_5945;
or2_5392: n_5938 <=  n_5939  OR n_5942;
and2_5393: n_5939 <=  n_5940  AND n_5941;
inv_5394: n_5940  <= TRANSPORT NOT a_N1120_aNOT_aOUT  ;
delay_5395: n_5941  <= TRANSPORT a_N1553_aQ  ;
and2_5396: n_5942 <=  n_5943  AND n_5944;
delay_5397: n_5943  <= TRANSPORT a_N130_aNOT_aOUT  ;
inv_5398: n_5944  <= TRANSPORT NOT a_N1120_aNOT_aOUT  ;
and1_5399: n_5945 <=  gnd;
delay_5400: a_LC5_A3_aOUT  <= TRANSPORT a_LC5_A3_aIN  ;
xor2_5401: a_LC5_A3_aIN <=  n_5948  XOR n_5955;
or2_5402: n_5948 <=  n_5949  OR n_5952;
and2_5403: n_5949 <=  n_5950  AND n_5951;
inv_5404: n_5950  <= TRANSPORT NOT a_N1117_aOUT  ;
delay_5405: n_5951  <= TRANSPORT a_N1556_aQ  ;
and2_5406: n_5952 <=  n_5953  AND n_5954;
delay_5407: n_5953  <= TRANSPORT a_LC4_A3_aOUT  ;
inv_5408: n_5954  <= TRANSPORT NOT a_N1556_aQ  ;
and1_5409: n_5955 <=  gnd;
delay_5410: a_LC1_A3_aOUT  <= TRANSPORT a_LC1_A3_aIN  ;
xor2_5411: a_LC1_A3_aIN <=  n_5958  XOR n_5968;
or3_5412: n_5958 <=  n_5959  OR n_5962  OR n_5965;
and2_5413: n_5959 <=  n_5960  AND n_5961;
inv_5414: n_5960  <= TRANSPORT NOT a_N1555_aQ  ;
delay_5415: n_5961  <= TRANSPORT a_LC5_A3_aOUT  ;
and2_5416: n_5962 <=  n_5963  AND n_5964;
delay_5417: n_5963  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5418: n_5964  <= TRANSPORT a_LC5_A3_aOUT  ;
and2_5419: n_5965 <=  n_5966  AND n_5967;
inv_5420: n_5966  <= TRANSPORT NOT a_N1120_aNOT_aOUT  ;
delay_5421: n_5967  <= TRANSPORT a_N1160_aOUT  ;
and1_5422: n_5968 <=  gnd;
delay_5423: a_LC5_A7_aOUT  <= TRANSPORT a_LC5_A7_aIN  ;
xor2_5424: a_LC5_A7_aIN <=  n_5971  XOR n_5977;
or1_5425: n_5971 <=  n_5972;
and4_5426: n_5972 <=  n_5973  AND n_5974  AND n_5975  AND n_5976;
inv_5427: n_5973  <= TRANSPORT NOT a_N132_aOUT  ;
delay_5428: n_5974  <= TRANSPORT a_N1194_aNOT_aOUT  ;
delay_5429: n_5975  <= TRANSPORT a_N1555_aQ  ;
inv_5430: n_5976  <= TRANSPORT NOT a_N1556_aQ  ;
and1_5431: n_5977 <=  gnd;
dff_5432: DFF_a8251
    PORT MAP ( D => a_N1556_aD, CLK => a_N1556_aCLK, CLRN => a_N1556_aCLRN,
          PRN => vcc, Q => a_N1556_aQ);
delay_5433: a_N1556_aCLRN  <= TRANSPORT nRESET  ;
xor2_5434: a_N1556_aD <=  n_5984  XOR n_5993;
or3_5435: n_5984 <=  n_5985  OR n_5987  OR n_5990;
and1_5436: n_5985 <=  n_5986;
delay_5437: n_5986  <= TRANSPORT a_N264_aNOT_aOUT  ;
and2_5438: n_5987 <=  n_5988  AND n_5989;
delay_5439: n_5988  <= TRANSPORT a_N1187_aOUT  ;
delay_5440: n_5989  <= TRANSPORT a_LC1_A3_aOUT  ;
and2_5441: n_5990 <=  n_5991  AND n_5992;
delay_5442: n_5991  <= TRANSPORT a_N1187_aOUT  ;
delay_5443: n_5992  <= TRANSPORT a_LC5_A7_aOUT  ;
and1_5444: n_5993 <=  gnd;
delay_5445: n_5994  <= TRANSPORT nRXC  ;
filter_5446: FILTER_a8251
    PORT MAP (IN1 => n_5994, Y => a_N1556_aCLK);
delay_5447: a_LC6_D13_aOUT  <= TRANSPORT a_LC6_D13_aIN  ;
xor2_5448: a_LC6_D13_aIN <=  n_5998  XOR n_6003;
or1_5449: n_5998 <=  n_5999;
and3_5450: n_5999 <=  n_6000  AND n_6001  AND n_6002;
inv_5451: n_6000  <= TRANSPORT NOT a_N1152_aNOT_aOUT  ;
delay_5452: n_6001  <= TRANSPORT a_N62_aQ  ;
delay_5453: n_6002  <= TRANSPORT a_N63_aQ  ;
and1_5454: n_6003 <=  gnd;
delay_5455: a_N108_aNOT_aOUT  <= TRANSPORT a_N108_aNOT_aIN  ;
xor2_5456: a_N108_aNOT_aIN <=  n_6006  XOR n_6013;
or2_5457: n_6006 <=  n_6007  OR n_6011;
and3_5458: n_6007 <=  n_6008  AND n_6009  AND n_6010;
delay_5459: n_6008  <= TRANSPORT a_N95_aNOT_aOUT  ;
inv_5460: n_6009  <= TRANSPORT NOT a_N1152_aNOT_aOUT  ;
delay_5461: n_6010  <= TRANSPORT a_N1146_aOUT  ;
and1_5462: n_6011 <=  n_6012;
inv_5463: n_6012  <= TRANSPORT NOT a_N87_aNOT_aOUT  ;
and1_5464: n_6013 <=  gnd;
delay_5465: mode_cmplt_aOUT  <= TRANSPORT mode_cmplt_aIN  ;
xor2_5466: mode_cmplt_aIN <=  n_6015  XOR n_6021;
or1_5467: n_6015 <=  n_6016;
and4_5468: n_6016 <=  n_6017  AND n_6018  AND n_6019  AND n_6020;
delay_5469: n_6017  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5470: n_6018  <= TRANSPORT a_N1754_aQ  ;
inv_5471: n_6019  <= TRANSPORT NOT a_N1757_aQ  ;
inv_5472: n_6020  <= TRANSPORT NOT a_N1756_aQ  ;
and1_5473: n_6021 <=  gnd;
delay_5474: a_LC6_D11_aOUT  <= TRANSPORT a_LC6_D11_aIN  ;
xor2_5475: a_LC6_D11_aIN <=  n_6025  XOR n_6034;
or2_5476: n_6025 <=  n_6026  OR n_6030;
and3_5477: n_6026 <=  n_6027  AND n_6028  AND n_6029;
delay_5478: n_6027  <= TRANSPORT a_N64_aQ  ;
inv_5479: n_6028  <= TRANSPORT NOT a_N61_aQ  ;
inv_5480: n_6029  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and3_5481: n_6030 <=  n_6031  AND n_6032  AND n_6033;
inv_5482: n_6031  <= TRANSPORT NOT EXTSYNCD  ;
delay_5483: n_6032  <= TRANSPORT a_N64_aQ  ;
inv_5484: n_6033  <= TRANSPORT NOT a_N61_aQ  ;
and1_5485: n_6034 <=  gnd;
delay_5486: a_LC5_D11_aOUT  <= TRANSPORT a_LC5_D11_aIN  ;
xor2_5487: a_LC5_D11_aIN <=  n_6037  XOR n_6045;
or2_5488: n_6037 <=  n_6038  OR n_6042;
and3_5489: n_6038 <=  n_6039  AND n_6040  AND n_6041;
delay_5490: n_6039  <= TRANSPORT a_N127_aOUT  ;
inv_5491: n_6040  <= TRANSPORT NOT a_N59_aQ  ;
delay_5492: n_6041  <= TRANSPORT mode_cmplt_aOUT  ;
and2_5493: n_6042 <=  n_6043  AND n_6044;
inv_5494: n_6043  <= TRANSPORT NOT a_N59_aQ  ;
delay_5495: n_6044  <= TRANSPORT a_LC6_D11_aOUT  ;
and1_5496: n_6045 <=  gnd;
delay_5497: a_LC7_D11_aOUT  <= TRANSPORT a_LC7_D11_aIN  ;
xor2_5498: a_LC7_D11_aIN <=  n_6048  XOR n_6056;
or3_5499: n_6048 <=  n_6049  OR n_6051  OR n_6054;
and1_5500: n_6049 <=  n_6050;
delay_5501: n_6050  <= TRANSPORT a_LC5_D11_aOUT  ;
and2_5502: n_6051 <=  n_6052  AND n_6053;
delay_5503: n_6052  <= TRANSPORT a_N1144_aNOT_aOUT  ;
inv_5504: n_6053  <= TRANSPORT NOT a_N1152_aNOT_aOUT  ;
and1_5505: n_6054 <=  n_6055;
delay_5506: n_6055  <= TRANSPORT a_N1164_aOUT  ;
and1_5507: n_6056 <=  gnd;
delay_5508: a_LC7_D10_aOUT  <= TRANSPORT a_LC7_D10_aIN  ;
xor2_5509: a_LC7_D10_aIN <=  n_6059  XOR n_6066;
or2_5510: n_6059 <=  n_6060  OR n_6062;
and1_5511: n_6060 <=  n_6061;
delay_5512: n_6061  <= TRANSPORT a_N108_aNOT_aOUT  ;
and3_5513: n_6062 <=  n_6063  AND n_6064  AND n_6065;
delay_5514: n_6063  <= TRANSPORT a_LC7_D11_aOUT  ;
inv_5515: n_6064  <= TRANSPORT NOT a_N62_aQ  ;
inv_5516: n_6065  <= TRANSPORT NOT a_N63_aQ  ;
and1_5517: n_6066 <=  gnd;
delay_5518: a_LC4_D8_aOUT  <= TRANSPORT a_LC4_D8_aIN  ;
xor2_5519: a_LC4_D8_aIN <=  n_6069  XOR n_6078;
or2_5520: n_6069 <=  n_6070  OR n_6074;
and3_5521: n_6070 <=  n_6071  AND n_6072  AND n_6073;
inv_5522: n_6071  <= TRANSPORT NOT a_N1149_aNOT_aOUT  ;
inv_5523: n_6072  <= TRANSPORT NOT a_N1163_aNOT_aOUT  ;
delay_5524: n_6073  <= TRANSPORT RXD  ;
and3_5525: n_6074 <=  n_6075  AND n_6076  AND n_6077;
inv_5526: n_6075  <= TRANSPORT NOT a_N1149_aNOT_aOUT  ;
inv_5527: n_6076  <= TRANSPORT NOT a_N1163_aNOT_aOUT  ;
inv_5528: n_6077  <= TRANSPORT NOT a_N751_aNOT_aOUT  ;
and1_5529: n_6078 <=  gnd;
delay_5530: a_N1158_aOUT  <= TRANSPORT a_N1158_aIN  ;
xor2_5531: a_N1158_aIN <=  n_6081  XOR n_6085;
or1_5532: n_6081 <=  n_6082;
and2_5533: n_6082 <=  n_6083  AND n_6084;
delay_5534: n_6083  <= TRANSPORT a_SMODE_OUT_F0_G_aQ  ;
inv_5535: n_6084  <= TRANSPORT NOT a_SMODE_OUT_F1_G_aQ  ;
and1_5536: n_6085 <=  gnd;
delay_5537: a_N745_aNOT_aOUT  <= TRANSPORT a_N745_aNOT_aIN  ;
xor2_5538: a_N745_aNOT_aIN <=  n_6088  XOR n_6098;
or3_5539: n_6088 <=  n_6089  OR n_6092  OR n_6095;
and2_5540: n_6089 <=  n_6090  AND n_6091;
inv_5541: n_6090  <= TRANSPORT NOT a_N735_aNOT_aOUT  ;
delay_5542: n_6091  <= TRANSPORT a_N1158_aOUT  ;
and2_5543: n_6092 <=  n_6093  AND n_6094;
inv_5544: n_6093  <= TRANSPORT NOT a_N735_aNOT_aOUT  ;
inv_5545: n_6094  <= TRANSPORT NOT a_SCMND_OUT_F2_G_aQ  ;
and2_5546: n_6095 <=  n_6096  AND n_6097;
inv_5547: n_6096  <= TRANSPORT NOT a_N735_aNOT_aOUT  ;
delay_5548: n_6097  <= TRANSPORT RXD  ;
and1_5549: n_6098 <=  gnd;
delay_5550: a_LC3_D8_aOUT  <= TRANSPORT a_LC3_D8_aIN  ;
xor2_5551: a_LC3_D8_aIN <=  n_6101  XOR n_6110;
or4_5552: n_6101 <=  n_6102  OR n_6104  OR n_6106  OR n_6108;
and1_5553: n_6102 <=  n_6103;
delay_5554: n_6103  <= TRANSPORT a_LC4_D8_aOUT  ;
and1_5555: n_6104 <=  n_6105;
delay_5556: n_6105  <= TRANSPORT a_N745_aNOT_aOUT  ;
and1_5557: n_6106 <=  n_6107;
inv_5558: n_6107  <= TRANSPORT NOT a_N89_aNOT_aOUT  ;
and1_5559: n_6108 <=  n_6109;
delay_5560: n_6109  <= TRANSPORT a_LC8_D21_aOUT  ;
and1_5561: n_6110 <=  gnd;
delay_5562: a_LC7_D7_aOUT  <= TRANSPORT a_LC7_D7_aIN  ;
xor2_5563: a_LC7_D7_aIN <=  n_6113  XOR n_6118;
or1_5564: n_6113 <=  n_6114;
and3_5565: n_6114 <=  n_6115  AND n_6116  AND n_6117;
inv_5566: n_6115  <= TRANSPORT NOT a_N1175_aNOT_aOUT  ;
inv_5567: n_6116  <= TRANSPORT NOT a_N61_aQ  ;
delay_5568: n_6117  <= TRANSPORT a_N63_aQ  ;
and1_5569: n_6118 <=  gnd;
delay_5570: a_N141_aNOT_aOUT  <= TRANSPORT a_N141_aNOT_aIN  ;
xor2_5571: a_N141_aNOT_aIN <=  n_6120  XOR n_6126;
or1_5572: n_6120 <=  n_6121;
and4_5573: n_6121 <=  n_6122  AND n_6123  AND n_6124  AND n_6125;
inv_5574: n_6122  <= TRANSPORT NOT a_N64_aQ  ;
delay_5575: n_6123  <= TRANSPORT a_N62_aQ  ;
delay_5576: n_6124  <= TRANSPORT a_N61_aQ  ;
inv_5577: n_6125  <= TRANSPORT NOT a_N63_aQ  ;
and1_5578: n_6126 <=  gnd;
delay_5579: a_N106_aNOT_aOUT  <= TRANSPORT a_N106_aNOT_aIN  ;
xor2_5580: a_N106_aNOT_aIN <=  n_6129  XOR n_6137;
or3_5581: n_6129 <=  n_6130  OR n_6133  OR n_6135;
and2_5582: n_6130 <=  n_6131  AND n_6132;
delay_5583: n_6131  <= TRANSPORT a_N95_aNOT_aOUT  ;
delay_5584: n_6132  <= TRANSPORT a_LC7_D7_aOUT  ;
and1_5585: n_6133 <=  n_6134;
delay_5586: n_6134  <= TRANSPORT a_N141_aNOT_aOUT  ;
and1_5587: n_6135 <=  n_6136;
delay_5588: n_6136  <= TRANSPORT a_N113_aNOT_aOUT  ;
and1_5589: n_6137 <=  gnd;
delay_5590: a_LC4_D10_aOUT  <= TRANSPORT a_LC4_D10_aIN  ;
xor2_5591: a_LC4_D10_aIN <=  n_6140  XOR n_6149;
or4_5592: n_6140 <=  n_6141  OR n_6143  OR n_6145  OR n_6147;
and1_5593: n_6141 <=  n_6142;
delay_5594: n_6142  <= TRANSPORT a_LC7_D10_aOUT  ;
and1_5595: n_6143 <=  n_6144;
delay_5596: n_6144  <= TRANSPORT a_LC3_D8_aOUT  ;
and1_5597: n_6145 <=  n_6146;
delay_5598: n_6146  <= TRANSPORT a_N106_aNOT_aOUT  ;
and1_5599: n_6147 <=  n_6148;
delay_5600: n_6148  <= TRANSPORT a_N743_aNOT_aOUT  ;
and1_5601: n_6149 <=  gnd;
delay_5602: a_LC5_D13_aOUT  <= TRANSPORT a_LC5_D13_aIN  ;
xor2_5603: a_LC5_D13_aIN <=  n_6152  XOR n_6161;
or3_5604: n_6152 <=  n_6153  OR n_6156  OR n_6159;
and2_5605: n_6153 <=  n_6154  AND n_6155;
delay_5606: n_6154  <= TRANSPORT a_LC6_D13_aOUT  ;
inv_5607: n_6155  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_5608: n_6156 <=  n_6157  AND n_6158;
delay_5609: n_6157  <= TRANSPORT a_N132_aOUT  ;
delay_5610: n_6158  <= TRANSPORT a_LC6_D13_aOUT  ;
and1_5611: n_6159 <=  n_6160;
delay_5612: n_6160  <= TRANSPORT a_LC4_D10_aOUT  ;
and1_5613: n_6161 <=  gnd;
delay_5614: a_N740_aNOT_aOUT  <= TRANSPORT a_N740_aNOT_aIN  ;
xor2_5615: a_N740_aNOT_aIN <=  n_6164  XOR n_6169;
or1_5616: n_6164 <=  n_6165;
and3_5617: n_6165 <=  n_6166  AND n_6167  AND n_6168;
delay_5618: n_6166  <= TRANSPORT a_N1120_aNOT_aOUT  ;
inv_5619: n_6167  <= TRANSPORT NOT a_N132_aOUT  ;
delay_5620: n_6168  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_5621: n_6169 <=  gnd;
dff_5622: DFF_a8251
    PORT MAP ( D => a_N64_aD, CLK => a_N64_aCLK, CLRN => a_N64_aCLRN, PRN => vcc,
          Q => a_N64_aQ);
delay_5623: a_N64_aCLRN  <= TRANSPORT nRESET  ;
xor2_5624: a_N64_aD <=  n_6176  XOR n_6184;
or2_5625: n_6176 <=  n_6177  OR n_6180;
and2_5626: n_6177 <=  n_6178  AND n_6179;
inv_5627: n_6178  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5628: n_6179  <= TRANSPORT a_LC5_D13_aOUT  ;
and3_5629: n_6180 <=  n_6181  AND n_6182  AND n_6183;
inv_5630: n_6181  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5631: n_6182  <= TRANSPORT NOT a_LC1_D2_aNOT_aOUT  ;
inv_5632: n_6183  <= TRANSPORT NOT a_N740_aNOT_aOUT  ;
and1_5633: n_6184 <=  gnd;
delay_5634: n_6185  <= TRANSPORT nRXC  ;
filter_5635: FILTER_a8251
    PORT MAP (IN1 => n_6185, Y => a_N64_aCLK);
dff_5636: DFF_a8251
    PORT MAP ( D => a_N1301_aD, CLK => a_N1301_aCLK, CLRN => a_N1301_aCLRN,
          PRN => vcc, Q => a_N1301_aQ);
delay_5637: a_N1301_aCLRN  <= TRANSPORT nRESET  ;
xor2_5638: a_N1301_aD <=  n_6193  XOR n_6202;
or2_5639: n_6193 <=  n_6194  OR n_6198;
and3_5640: n_6194 <=  n_6195  AND n_6196  AND n_6197;
inv_5641: n_6195  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5642: n_6196  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5643: n_6197  <= TRANSPORT a_N1300_aQ  ;
and3_5644: n_6198 <=  n_6199  AND n_6200  AND n_6201;
inv_5645: n_6199  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5646: n_6200  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5647: n_6201  <= TRANSPORT a_N1301_aQ  ;
and1_5648: n_6202 <=  gnd;
delay_5649: n_6203  <= TRANSPORT nRXC  ;
filter_5650: FILTER_a8251
    PORT MAP (IN1 => n_6203, Y => a_N1301_aCLK);
dff_5651: DFF_a8251
    PORT MAP ( D => a_N1998_aD, CLK => a_N1998_aCLK, CLRN => a_N1998_aCLRN,
          PRN => vcc, Q => a_N1998_aQ);
delay_5652: a_N1998_aCLRN  <= TRANSPORT nRESET  ;
xor2_5653: a_N1998_aD <=  n_6211  XOR n_6220;
or2_5654: n_6211 <=  n_6212  OR n_6216;
and3_5655: n_6212 <=  n_6213  AND n_6214  AND n_6215;
inv_5656: n_6213  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5657: n_6214  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5658: n_6215  <= TRANSPORT a_N1998_aQ  ;
and3_5659: n_6216 <=  n_6217  AND n_6218  AND n_6219;
inv_5660: n_6217  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5661: n_6218  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5662: n_6219  <= TRANSPORT RXD  ;
and1_5663: n_6220 <=  gnd;
delay_5664: n_6221  <= TRANSPORT nRXC  ;
filter_5665: FILTER_a8251
    PORT MAP (IN1 => n_6221, Y => a_N1998_aCLK);
dff_5666: DFF_a8251
    PORT MAP ( D => a_N1300_aD, CLK => a_N1300_aCLK, CLRN => a_N1300_aCLRN,
          PRN => vcc, Q => a_N1300_aQ);
delay_5667: a_N1300_aCLRN  <= TRANSPORT nRESET  ;
xor2_5668: a_N1300_aD <=  n_6229  XOR n_6238;
or2_5669: n_6229 <=  n_6230  OR n_6234;
and3_5670: n_6230 <=  n_6231  AND n_6232  AND n_6233;
inv_5671: n_6231  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5672: n_6232  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5673: n_6233  <= TRANSPORT a_N1998_aQ  ;
and3_5674: n_6234 <=  n_6235  AND n_6236  AND n_6237;
inv_5675: n_6235  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5676: n_6236  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5677: n_6237  <= TRANSPORT a_N1300_aQ  ;
and1_5678: n_6238 <=  gnd;
delay_5679: n_6239  <= TRANSPORT nRXC  ;
filter_5680: FILTER_a8251
    PORT MAP (IN1 => n_6239, Y => a_N1300_aCLK);
dff_5681: DFF_a8251
    PORT MAP ( D => a_N2031_aD, CLK => a_N2031_aCLK, CLRN => a_N2031_aCLRN,
          PRN => vcc, Q => a_N2031_aQ);
delay_5682: a_N2031_aCLRN  <= TRANSPORT nRESET  ;
xor2_5683: a_N2031_aD <=  n_6247  XOR n_6254;
or2_5684: n_6247 <=  n_6248  OR n_6251;
and2_5685: n_6248 <=  n_6249  AND n_6250;
delay_5686: n_6249  <= TRANSPORT a_N1197_aOUT  ;
delay_5687: n_6250  <= TRANSPORT DIN(0)  ;
and2_5688: n_6251 <=  n_6252  AND n_6253;
delay_5689: n_6252  <= TRANSPORT a_N1198_aOUT  ;
delay_5690: n_6253  <= TRANSPORT a_N2031_aQ  ;
and1_5691: n_6254 <=  gnd;
inv_5692: n_6255  <= TRANSPORT NOT nTXC  ;
filter_5693: FILTER_a8251
    PORT MAP (IN1 => n_6255, Y => a_N2031_aCLK);
delay_5694: a_N1123_aNOT_aOUT  <= TRANSPORT a_N1123_aNOT_aIN  ;
xor2_5695: a_N1123_aNOT_aIN <=  n_6258  XOR n_6265;
or3_5696: n_6258 <=  n_6259  OR n_6261  OR n_6263;
and1_5697: n_6259 <=  n_6260;
delay_5698: n_6260  <= TRANSPORT a_N1756_aQ  ;
and1_5699: n_6261 <=  n_6262;
delay_5700: n_6262  <= TRANSPORT a_N1757_aQ  ;
and1_5701: n_6263 <=  n_6264;
delay_5702: n_6264  <= TRANSPORT a_N1754_aQ  ;
and1_5703: n_6265 <=  gnd;
delay_5704: a_LC3_C8_aOUT  <= TRANSPORT a_LC3_C8_aIN  ;
xor2_5705: a_LC3_C8_aIN <=  n_6268  XOR n_6274;
or1_5706: n_6268 <=  n_6269;
and4_5707: n_6269 <=  n_6270  AND n_6271  AND n_6272  AND n_6273;
delay_5708: n_6270  <= TRANSPORT a_N1189_aOUT  ;
delay_5709: n_6271  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_5710: n_6272  <= TRANSPORT NOT a_N1123_aNOT_aOUT  ;
delay_5711: n_6273  <= TRANSPORT DIN(5)  ;
and1_5712: n_6274 <=  gnd;
delay_5713: a_N1034_aNOT_aOUT  <= TRANSPORT a_N1034_aNOT_aIN  ;
xor2_5714: a_N1034_aNOT_aIN <=  n_6276  XOR n_6283;
or3_5715: n_6276 <=  n_6277  OR n_6279  OR n_6281;
and1_5716: n_6277 <=  n_6278;
delay_5717: n_6278  <= TRANSPORT a_N1123_aNOT_aOUT  ;
and1_5718: n_6279 <=  n_6280;
inv_5719: n_6280  <= TRANSPORT NOT a_N82_aNOT_aOUT  ;
and1_5720: n_6281 <=  n_6282;
inv_5721: n_6282  <= TRANSPORT NOT a_N1189_aOUT  ;
and1_5722: n_6283 <=  gnd;
dff_5723: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F5_G_aD, CLK => a_SMODE_OUT_F5_G_aCLK, CLRN => a_SMODE_OUT_F5_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F5_G_aQ);
delay_5724: a_SMODE_OUT_F5_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_5725: a_SMODE_OUT_F5_G_aD <=  n_6290  XOR n_6298;
or2_5726: n_6290 <=  n_6291  OR n_6294;
and2_5727: n_6291 <=  n_6292  AND n_6293;
delay_5728: n_6292  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5729: n_6293  <= TRANSPORT a_LC3_C8_aOUT  ;
and3_5730: n_6294 <=  n_6295  AND n_6296  AND n_6297;
delay_5731: n_6295  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5732: n_6296  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_5733: n_6297  <= TRANSPORT a_SMODE_OUT_F5_G_aQ  ;
and1_5734: n_6298 <=  gnd;
delay_5735: n_6299  <= TRANSPORT CLK  ;
filter_5736: FILTER_a8251
    PORT MAP (IN1 => n_6299, Y => a_SMODE_OUT_F5_G_aCLK);
delay_5737: a_N317_aOUT  <= TRANSPORT a_N317_aIN  ;
xor2_5738: a_N317_aIN <=  n_6303  XOR n_6307;
or1_5739: n_6303 <=  n_6304;
and2_5740: n_6304 <=  n_6305  AND n_6306;
inv_5741: n_6305  <= TRANSPORT NOT a_N470_aOUT  ;
delay_5742: n_6306  <= TRANSPORT a_N397_aQ  ;
and1_5743: n_6307 <=  gnd;
dff_5744: DFF_a8251
    PORT MAP ( D => a_N394_aD, CLK => a_N394_aCLK, CLRN => a_N394_aCLRN, PRN => vcc,
          Q => a_N394_aQ);
delay_5745: a_N394_aCLRN  <= TRANSPORT nRESET  ;
xor2_5746: a_N394_aD <=  n_6314  XOR n_6328;
or3_5747: n_6314 <=  n_6315  OR n_6319  OR n_6323;
and3_5748: n_6315 <=  n_6316  AND n_6317  AND n_6318;
delay_5749: n_6316  <= TRANSPORT a_N1056_aOUT  ;
inv_5750: n_6317  <= TRANSPORT NOT a_N317_aOUT  ;
delay_5751: n_6318  <= TRANSPORT a_N394_aQ  ;
and3_5752: n_6319 <=  n_6320  AND n_6321  AND n_6322;
delay_5753: n_6320  <= TRANSPORT a_N1056_aOUT  ;
inv_5754: n_6321  <= TRANSPORT NOT a_N396_aQ  ;
delay_5755: n_6322  <= TRANSPORT a_N394_aQ  ;
and4_5756: n_6323 <=  n_6324  AND n_6325  AND n_6326  AND n_6327;
delay_5757: n_6324  <= TRANSPORT a_N1056_aOUT  ;
delay_5758: n_6325  <= TRANSPORT a_N396_aQ  ;
delay_5759: n_6326  <= TRANSPORT a_N317_aOUT  ;
inv_5760: n_6327  <= TRANSPORT NOT a_N394_aQ  ;
and1_5761: n_6328 <=  gnd;
inv_5762: n_6329  <= TRANSPORT NOT nTXC  ;
filter_5763: FILTER_a8251
    PORT MAP (IN1 => n_6329, Y => a_N394_aCLK);
delay_5764: a_N1067_aOUT  <= TRANSPORT a_N1067_aIN  ;
xor2_5765: a_N1067_aIN <=  n_6333  XOR n_6339;
or1_5766: n_6333 <=  n_6334;
and4_5767: n_6334 <=  n_6335  AND n_6336  AND n_6337  AND n_6338;
inv_5768: n_6335  <= TRANSPORT NOT a_N1175_aNOT_aOUT  ;
delay_5769: n_6336  <= TRANSPORT a_N132_aOUT  ;
delay_5770: n_6337  <= TRANSPORT a_N61_aQ  ;
delay_5771: n_6338  <= TRANSPORT a_N63_aQ  ;
and1_5772: n_6339 <=  gnd;
delay_5773: a_LC3_D10_aOUT  <= TRANSPORT a_LC3_D10_aIN  ;
xor2_5774: a_LC3_D10_aIN <=  n_6342  XOR n_6351;
or4_5775: n_6342 <=  n_6343  OR n_6345  OR n_6347  OR n_6349;
and1_5776: n_6343 <=  n_6344;
delay_5777: n_6344  <= TRANSPORT a_N106_aNOT_aOUT  ;
and1_5778: n_6345 <=  n_6346;
inv_5779: n_6346  <= TRANSPORT NOT a_N247_aNOT_aOUT  ;
and1_5780: n_6347 <=  n_6348;
inv_5781: n_6348  <= TRANSPORT NOT a_LC1_D14_aNOT_aOUT  ;
and1_5782: n_6349 <=  n_6350;
inv_5783: n_6350  <= TRANSPORT NOT a_N1073_aNOT_aOUT  ;
and1_5784: n_6351 <=  gnd;
delay_5785: a_LC2_D13_aOUT  <= TRANSPORT a_LC2_D13_aIN  ;
xor2_5786: a_LC2_D13_aIN <=  n_6354  XOR n_6362;
or3_5787: n_6354 <=  n_6355  OR n_6357  OR n_6360;
and1_5788: n_6355 <=  n_6356;
delay_5789: n_6356  <= TRANSPORT a_N1067_aOUT  ;
and2_5790: n_6357 <=  n_6358  AND n_6359;
delay_5791: n_6358  <= TRANSPORT a_N132_aOUT  ;
delay_5792: n_6359  <= TRANSPORT a_N1080_aOUT  ;
and1_5793: n_6360 <=  n_6361;
delay_5794: n_6361  <= TRANSPORT a_LC3_D10_aOUT  ;
and1_5795: n_6362 <=  gnd;
delay_5796: a_LC4_D13_aOUT  <= TRANSPORT a_LC4_D13_aIN  ;
xor2_5797: a_LC4_D13_aIN <=  n_6365  XOR n_6373;
or2_5798: n_6365 <=  n_6366  OR n_6369;
and2_5799: n_6366 <=  n_6367  AND n_6368;
inv_5800: n_6367  <= TRANSPORT NOT a_N64_aQ  ;
delay_5801: n_6368  <= TRANSPORT a_N62_aQ  ;
and3_5802: n_6369 <=  n_6370  AND n_6371  AND n_6372;
delay_5803: n_6370  <= TRANSPORT a_N740_aNOT_aOUT  ;
delay_5804: n_6371  <= TRANSPORT a_N64_aQ  ;
inv_5805: n_6372  <= TRANSPORT NOT a_N62_aQ  ;
and1_5806: n_6373 <=  gnd;
dff_5807: DFF_a8251
    PORT MAP ( D => a_N62_aD, CLK => a_N62_aCLK, CLRN => a_N62_aCLRN, PRN => vcc,
          Q => a_N62_aQ);
delay_5808: a_N62_aCLRN  <= TRANSPORT nRESET  ;
xor2_5809: a_N62_aD <=  n_6380  XOR n_6388;
or2_5810: n_6380 <=  n_6381  OR n_6384;
and2_5811: n_6381 <=  n_6382  AND n_6383;
inv_5812: n_6382  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5813: n_6383  <= TRANSPORT a_LC2_D13_aOUT  ;
and3_5814: n_6384 <=  n_6385  AND n_6386  AND n_6387;
inv_5815: n_6385  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5816: n_6386  <= TRANSPORT NOT a_N1118_aNOT_aOUT  ;
delay_5817: n_6387  <= TRANSPORT a_LC4_D13_aOUT  ;
and1_5818: n_6388 <=  gnd;
delay_5819: n_6389  <= TRANSPORT nRXC  ;
filter_5820: FILTER_a8251
    PORT MAP (IN1 => n_6389, Y => a_N62_aCLK);
delay_5821: a_LC1_C7_aNOT_aOUT  <= TRANSPORT a_LC1_C7_aNOT_aIN  ;
xor2_5822: a_LC1_C7_aNOT_aIN <=  n_6392  XOR n_6397;
or1_5823: n_6392 <=  n_6393;
and3_5824: n_6393 <=  n_6394  AND n_6395  AND n_6396;
delay_5825: n_6394  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5826: n_6395  <= TRANSPORT a_N1806_aQ  ;
inv_5827: n_6396  <= TRANSPORT NOT a_N1808_aQ  ;
and1_5828: n_6397 <=  gnd;
delay_5829: a_N1121_aNOT_aOUT  <= TRANSPORT a_N1121_aNOT_aIN  ;
xor2_5830: a_N1121_aNOT_aIN <=  n_6399  XOR n_6405;
or2_5831: n_6399 <=  n_6400  OR n_6403;
and2_5832: n_6400 <=  n_6401  AND n_6402;
delay_5833: n_6401  <= TRANSPORT a_N1898_aQ  ;
inv_5834: n_6402  <= TRANSPORT NOT a_N1897_aQ  ;
and1_5835: n_6403 <=  n_6404;
delay_5836: n_6404  <= TRANSPORT a_N83_aOUT  ;
and1_5837: n_6405 <=  gnd;
delay_5838: a_N701_aNOT_aOUT  <= TRANSPORT a_N701_aNOT_aIN  ;
xor2_5839: a_N701_aNOT_aIN <=  n_6407  XOR n_6411;
or1_5840: n_6407 <=  n_6408;
and2_5841: n_6408 <=  n_6409  AND n_6410;
delay_5842: n_6409  <= TRANSPORT a_LC1_C7_aNOT_aOUT  ;
inv_5843: n_6410  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
and1_5844: n_6411 <=  gnd;
delay_5845: a_N611_aOUT  <= TRANSPORT a_N611_aIN  ;
xor2_5846: a_N611_aIN <=  n_6414  XOR n_6418;
or1_5847: n_6414 <=  n_6415;
and2_5848: n_6415 <=  n_6416  AND n_6417;
delay_5849: n_6416  <= TRANSPORT DIN(7)  ;
delay_5850: n_6417  <= TRANSPORT a_N701_aNOT_aOUT  ;
and1_5851: n_6418 <=  gnd;
delay_5852: a_N613_aOUT  <= TRANSPORT a_N613_aIN  ;
xor2_5853: a_N613_aIN <=  n_6420  XOR n_6429;
or3_5854: n_6420 <=  n_6421  OR n_6423  OR n_6426;
and1_5855: n_6421 <=  n_6422;
delay_5856: n_6422  <= TRANSPORT a_N1121_aNOT_aOUT  ;
and2_5857: n_6423 <=  n_6424  AND n_6425;
delay_5858: n_6424  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_5859: n_6425  <= TRANSPORT a_N1808_aQ  ;
and2_5860: n_6426 <=  n_6427  AND n_6428;
delay_5861: n_6427  <= TRANSPORT a_N1120_aNOT_aOUT  ;
inv_5862: n_6428  <= TRANSPORT NOT a_N1806_aQ  ;
and1_5863: n_6429 <=  gnd;
dff_5864: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F7_G_aD, CLK => a_SCMND_OUT_F7_G_aCLK, CLRN => a_SCMND_OUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F7_G_aQ);
delay_5865: a_SCMND_OUT_F7_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_5866: a_SCMND_OUT_F7_G_aD <=  n_6437  XOR n_6445;
or2_5867: n_6437 <=  n_6438  OR n_6441;
and2_5868: n_6438 <=  n_6439  AND n_6440;
delay_5869: n_6439  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5870: n_6440  <= TRANSPORT a_N611_aOUT  ;
and3_5871: n_6441 <=  n_6442  AND n_6443  AND n_6444;
delay_5872: n_6442  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5873: n_6443  <= TRANSPORT a_N613_aOUT  ;
delay_5874: n_6444  <= TRANSPORT a_SCMND_OUT_F7_G_aQ  ;
and1_5875: n_6445 <=  gnd;
delay_5876: n_6446  <= TRANSPORT CLK  ;
filter_5877: FILTER_a8251
    PORT MAP (IN1 => n_6446, Y => a_SCMND_OUT_F7_G_aCLK);
dff_5878: DFF_a8251
    PORT MAP ( D => a_N1902_aD, CLK => a_N1902_aCLK, CLRN => a_N1902_aCLRN,
          PRN => vcc, Q => a_N1902_aQ);
delay_5879: a_N1902_aCLRN  <= TRANSPORT nRESET  ;
xor2_5880: a_N1902_aD <=  n_6454  XOR n_6457;
or1_5881: n_6454 <=  n_6455;
and1_5882: n_6455 <=  n_6456;
delay_5883: n_6456  <= TRANSPORT a_N1902_aQ  ;
and1_5884: n_6457 <=  gnd;
delay_5885: n_6458  <= TRANSPORT nRXC  ;
filter_5886: FILTER_a8251
    PORT MAP (IN1 => n_6458, Y => a_N1902_aCLK);
dff_5887: DFF_a8251
    PORT MAP ( D => a_N1901_aD, CLK => a_N1901_aCLK, CLRN => a_N1901_aCLRN,
          PRN => vcc, Q => a_N1901_aQ);
delay_5888: a_N1901_aCLRN  <= TRANSPORT nRESET  ;
xor2_5889: a_N1901_aD <=  n_6466  XOR n_6469;
or1_5890: n_6466 <=  n_6467;
and1_5891: n_6467 <=  n_6468;
delay_5892: n_6468  <= TRANSPORT a_SCMND_OUT_F7_G_aQ  ;
and1_5893: n_6469 <=  gnd;
delay_5894: n_6470  <= TRANSPORT nRXC  ;
filter_5895: FILTER_a8251
    PORT MAP (IN1 => n_6470, Y => a_N1901_aCLK);
dff_5896: DFF_a8251
    PORT MAP ( D => a_N1305_aD, CLK => a_N1305_aCLK, CLRN => a_N1305_aCLRN,
          PRN => vcc, Q => a_N1305_aQ);
delay_5897: a_N1305_aCLRN  <= TRANSPORT nRESET  ;
xor2_5898: a_N1305_aD <=  n_6478  XOR n_6487;
or2_5899: n_6478 <=  n_6479  OR n_6483;
and3_5900: n_6479 <=  n_6480  AND n_6481  AND n_6482;
inv_5901: n_6480  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5902: n_6481  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5903: n_6482  <= TRANSPORT a_N1305_aQ  ;
and3_5904: n_6483 <=  n_6484  AND n_6485  AND n_6486;
inv_5905: n_6484  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5906: n_6485  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5907: n_6486  <= TRANSPORT a_N1304_aQ  ;
and1_5908: n_6487 <=  gnd;
delay_5909: n_6488  <= TRANSPORT nRXC  ;
filter_5910: FILTER_a8251
    PORT MAP (IN1 => n_6488, Y => a_N1305_aCLK);
dff_5911: DFF_a8251
    PORT MAP ( D => a_N1304_aD, CLK => a_N1304_aCLK, CLRN => a_N1304_aCLRN,
          PRN => vcc, Q => a_N1304_aQ);
delay_5912: a_N1304_aCLRN  <= TRANSPORT nRESET  ;
xor2_5913: a_N1304_aD <=  n_6496  XOR n_6505;
or2_5914: n_6496 <=  n_6497  OR n_6501;
and3_5915: n_6497 <=  n_6498  AND n_6499  AND n_6500;
inv_5916: n_6498  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5917: n_6499  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5918: n_6500  <= TRANSPORT a_N1303_aQ  ;
and3_5919: n_6501 <=  n_6502  AND n_6503  AND n_6504;
inv_5920: n_6502  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5921: n_6503  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5922: n_6504  <= TRANSPORT a_N1304_aQ  ;
and1_5923: n_6505 <=  gnd;
delay_5924: n_6506  <= TRANSPORT nRXC  ;
filter_5925: FILTER_a8251
    PORT MAP (IN1 => n_6506, Y => a_N1304_aCLK);
dff_5926: DFF_a8251
    PORT MAP ( D => a_N1303_aD, CLK => a_N1303_aCLK, CLRN => a_N1303_aCLRN,
          PRN => vcc, Q => a_N1303_aQ);
delay_5927: a_N1303_aCLRN  <= TRANSPORT nRESET  ;
xor2_5928: a_N1303_aD <=  n_6514  XOR n_6523;
or2_5929: n_6514 <=  n_6515  OR n_6519;
and3_5930: n_6515 <=  n_6516  AND n_6517  AND n_6518;
inv_5931: n_6516  <= TRANSPORT NOT a_N83_aOUT  ;
inv_5932: n_6517  <= TRANSPORT NOT a_N1124_aNOT_aOUT  ;
delay_5933: n_6518  <= TRANSPORT a_N1303_aQ  ;
and3_5934: n_6519 <=  n_6520  AND n_6521  AND n_6522;
inv_5935: n_6520  <= TRANSPORT NOT a_N83_aOUT  ;
delay_5936: n_6521  <= TRANSPORT a_N1124_aNOT_aOUT  ;
delay_5937: n_6522  <= TRANSPORT a_N1302_aQ  ;
and1_5938: n_6523 <=  gnd;
delay_5939: n_6524  <= TRANSPORT nRXC  ;
filter_5940: FILTER_a8251
    PORT MAP (IN1 => n_6524, Y => a_N1303_aCLK);
delay_5941: a_LC3_C3_aOUT  <= TRANSPORT a_LC3_C3_aIN  ;
xor2_5942: a_LC3_C3_aIN <=  n_6528  XOR n_6533;
or1_5943: n_6528 <=  n_6529;
and3_5944: n_6529 <=  n_6530  AND n_6531  AND n_6532;
delay_5945: n_6530  <= TRANSPORT a_N1189_aOUT  ;
delay_5946: n_6531  <= TRANSPORT DIN(7)  ;
inv_5947: n_6532  <= TRANSPORT NOT a_N1123_aNOT_aOUT  ;
and1_5948: n_6533 <=  gnd;
dff_5949: DFF_a8251
    PORT MAP ( D => a_SMODE_OUT_F7_G_aD, CLK => a_SMODE_OUT_F7_G_aCLK, CLRN => a_SMODE_OUT_F7_G_aCLRN,
          PRN => vcc, Q => a_SMODE_OUT_F7_G_aQ);
delay_5950: a_SMODE_OUT_F7_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_5951: a_SMODE_OUT_F7_G_aD <=  n_6540  XOR n_6548;
or2_5952: n_6540 <=  n_6541  OR n_6545;
and3_5953: n_6541 <=  n_6542  AND n_6543  AND n_6544;
delay_5954: n_6542  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5955: n_6543  <= TRANSPORT a_N1034_aNOT_aOUT  ;
delay_5956: n_6544  <= TRANSPORT a_SMODE_OUT_F7_G_aQ  ;
and2_5957: n_6545 <=  n_6546  AND n_6547;
delay_5958: n_6546  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_5959: n_6547  <= TRANSPORT a_LC3_C3_aOUT  ;
and1_5960: n_6548 <=  gnd;
delay_5961: n_6549  <= TRANSPORT CLK  ;
filter_5962: FILTER_a8251
    PORT MAP (IN1 => n_6549, Y => a_SMODE_OUT_F7_G_aCLK);
delay_5963: a_LC1_A8_aOUT  <= TRANSPORT a_LC1_A8_aIN  ;
xor2_5964: a_LC1_A8_aIN <=  n_6553  XOR n_6566;
or4_5965: n_6553 <=  n_6554  OR n_6557  OR n_6560  OR n_6563;
and1_5966: n_6554 <=  n_6555;
delay_5967: n_6555  <= TRANSPORT a_N965_aQ  ;
and1_5968: n_6557 <=  n_6558;
inv_5969: n_6558  <= TRANSPORT NOT a_N963_aQ  ;
and1_5970: n_6560 <=  n_6561;
inv_5971: n_6561  <= TRANSPORT NOT a_N964_aQ  ;
and1_5972: n_6563 <=  n_6564;
delay_5973: n_6564  <= TRANSPORT a_N962_aQ  ;
and1_5974: n_6566 <=  gnd;
delay_5975: a_LC4_A8_aOUT  <= TRANSPORT a_LC4_A8_aIN  ;
xor2_5976: a_LC4_A8_aIN <=  n_6569  XOR n_6579;
or3_5977: n_6569 <=  n_6570  OR n_6573  OR n_6576;
and2_5978: n_6570 <=  n_6571  AND n_6572;
inv_5979: n_6571  <= TRANSPORT NOT a_N1134_aNOT_aOUT  ;
inv_5980: n_6572  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_5981: n_6573 <=  n_6574  AND n_6575;
inv_5982: n_6574  <= TRANSPORT NOT a_N35_aNOT_aOUT  ;
inv_5983: n_6575  <= TRANSPORT NOT a_N963_aQ  ;
and2_5984: n_6576 <=  n_6577  AND n_6578;
delay_5985: n_6577  <= TRANSPORT a_N35_aNOT_aOUT  ;
delay_5986: n_6578  <= TRANSPORT a_N963_aQ  ;
and1_5987: n_6579 <=  gnd;
delay_5988: a_LC3_A8_aOUT  <= TRANSPORT a_LC3_A8_aIN  ;
xor2_5989: a_LC3_A8_aIN <=  n_6582  XOR n_6595;
or4_5990: n_6582 <=  n_6583  OR n_6585  OR n_6589  OR n_6592;
and1_5991: n_6583 <=  n_6584;
inv_5992: n_6584  <= TRANSPORT NOT a_N962_aQ  ;
and3_5993: n_6585 <=  n_6586  AND n_6587  AND n_6588;
delay_5994: n_6586  <= TRANSPORT a_N1134_aNOT_aOUT  ;
inv_5995: n_6587  <= TRANSPORT NOT a_N1052_aOUT  ;
delay_5996: n_6588  <= TRANSPORT a_N964_aQ  ;
and2_5997: n_6589 <=  n_6590  AND n_6591;
delay_5998: n_6590  <= TRANSPORT a_N1052_aOUT  ;
inv_5999: n_6591  <= TRANSPORT NOT a_N964_aQ  ;
and2_6000: n_6592 <=  n_6593  AND n_6594;
inv_6001: n_6593  <= TRANSPORT NOT a_N1134_aNOT_aOUT  ;
inv_6002: n_6594  <= TRANSPORT NOT a_N964_aQ  ;
and1_6003: n_6595 <=  gnd;
delay_6004: a_N383_aOUT  <= TRANSPORT a_N383_aIN  ;
xor2_6005: a_N383_aIN <=  n_6598  XOR n_6607;
or4_6006: n_6598 <=  n_6599  OR n_6601  OR n_6603  OR n_6605;
and1_6007: n_6599 <=  n_6600;
inv_6008: n_6600  <= TRANSPORT NOT a_N965_aQ  ;
and1_6009: n_6601 <=  n_6602;
inv_6010: n_6602  <= TRANSPORT NOT a_N964_aQ  ;
and1_6011: n_6603 <=  n_6604;
delay_6012: n_6604  <= TRANSPORT a_N962_aQ  ;
and1_6013: n_6605 <=  n_6606;
delay_6014: n_6606  <= TRANSPORT a_N35_aNOT_aOUT  ;
and1_6015: n_6607 <=  gnd;
delay_6016: a_LC2_A8_aOUT  <= TRANSPORT a_LC2_A8_aIN  ;
xor2_6017: a_LC2_A8_aIN <=  n_6610  XOR n_6630;
or5_6018: n_6610 <=  n_6611  OR n_6615  OR n_6619  OR n_6622  OR n_6626;
and3_6019: n_6611 <=  n_6612  AND n_6613  AND n_6614;
delay_6020: n_6612  <= TRANSPORT a_N965_aQ  ;
delay_6021: n_6613  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
delay_6022: n_6614  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and3_6023: n_6615 <=  n_6616  AND n_6617  AND n_6618;
delay_6024: n_6616  <= TRANSPORT a_N965_aQ  ;
inv_6025: n_6617  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
inv_6026: n_6618  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_6027: n_6619 <=  n_6620  AND n_6621;
delay_6028: n_6620  <= TRANSPORT a_N965_aQ  ;
inv_6029: n_6621  <= TRANSPORT NOT a_SMODE_OUT_F3_G_aQ  ;
and3_6030: n_6622 <=  n_6623  AND n_6624  AND n_6625;
inv_6031: n_6623  <= TRANSPORT NOT a_N965_aQ  ;
delay_6032: n_6624  <= TRANSPORT a_SMODE_OUT_F2_G_aQ  ;
inv_6033: n_6625  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and3_6034: n_6626 <=  n_6627  AND n_6628  AND n_6629;
inv_6035: n_6627  <= TRANSPORT NOT a_N965_aQ  ;
inv_6036: n_6628  <= TRANSPORT NOT a_SMODE_OUT_F2_G_aQ  ;
delay_6037: n_6629  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and1_6038: n_6630 <=  gnd;
delay_6039: a_N390_aOUT  <= TRANSPORT a_N390_aIN  ;
xor2_6040: a_N390_aIN <=  n_6633  XOR n_6642;
or3_6041: n_6633 <=  n_6634  OR n_6636  OR n_6639;
and1_6042: n_6634 <=  n_6635;
delay_6043: n_6635  <= TRANSPORT a_LC4_A8_aOUT  ;
and2_6044: n_6636 <=  n_6637  AND n_6638;
delay_6045: n_6637  <= TRANSPORT a_LC3_A8_aOUT  ;
delay_6046: n_6638  <= TRANSPORT a_N383_aOUT  ;
and2_6047: n_6639 <=  n_6640  AND n_6641;
delay_6048: n_6640  <= TRANSPORT a_N383_aOUT  ;
delay_6049: n_6641  <= TRANSPORT a_LC2_A8_aOUT  ;
and1_6050: n_6642 <=  gnd;
delay_6051: a_N143_aOUT  <= TRANSPORT a_N143_aIN  ;
xor2_6052: a_N143_aIN <=  n_6644  XOR n_6654;
or3_6053: n_6644 <=  n_6645  OR n_6648  OR n_6651;
and2_6054: n_6645 <=  n_6646  AND n_6647;
delay_6055: n_6646  <= TRANSPORT a_LC1_A8_aOUT  ;
delay_6056: n_6647  <= TRANSPORT a_N390_aOUT  ;
and2_6057: n_6648 <=  n_6649  AND n_6650;
delay_6058: n_6649  <= TRANSPORT a_N390_aOUT  ;
delay_6059: n_6650  <= TRANSPORT a_SMODE_OUT_F4_G_aQ  ;
and2_6060: n_6651 <=  n_6652  AND n_6653;
delay_6061: n_6652  <= TRANSPORT a_N1134_aNOT_aOUT  ;
delay_6062: n_6653  <= TRANSPORT a_N390_aOUT  ;
and1_6063: n_6654 <=  gnd;
delay_6064: a_LC1_A6_aOUT  <= TRANSPORT a_LC1_A6_aIN  ;
xor2_6065: a_LC1_A6_aIN <=  n_6657  XOR n_6661;
or1_6066: n_6657 <=  n_6658;
and2_6067: n_6658 <=  n_6659  AND n_6660;
inv_6068: n_6659  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_6069: n_6660  <= TRANSPORT RXD  ;
and1_6070: n_6661 <=  gnd;
delay_6071: a_N451_aOUT  <= TRANSPORT a_N451_aIN  ;
xor2_6072: a_N451_aIN <=  n_6664  XOR n_6671;
or2_6073: n_6664 <=  n_6665  OR n_6669;
and3_6074: n_6665 <=  n_6666  AND n_6667  AND n_6668;
inv_6075: n_6666  <= TRANSPORT NOT a_N129_aNOT_aOUT  ;
inv_6076: n_6667  <= TRANSPORT NOT a_LC8_A9_aOUT  ;
delay_6077: n_6668  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_6078: n_6669 <=  n_6670;
delay_6079: n_6670  <= TRANSPORT a_N1158_aOUT  ;
and1_6080: n_6671 <=  gnd;
dff_6081: DFF_a8251
    PORT MAP ( D => a_N965_aD, CLK => a_N965_aCLK, CLRN => a_N965_aCLRN, PRN => vcc,
          Q => a_N965_aQ);
delay_6082: a_N965_aCLRN  <= TRANSPORT nRESET  ;
xor2_6083: a_N965_aD <=  n_6678  XOR n_6692;
or3_6084: n_6678 <=  n_6679  OR n_6683  OR n_6687;
and3_6085: n_6679 <=  n_6680  AND n_6681  AND n_6682;
inv_6086: n_6680  <= TRANSPORT NOT a_N143_aOUT  ;
delay_6087: n_6681  <= TRANSPORT a_LC1_A6_aOUT  ;
delay_6088: n_6682  <= TRANSPORT a_N965_aQ  ;
and3_6089: n_6683 <=  n_6684  AND n_6685  AND n_6686;
delay_6090: n_6684  <= TRANSPORT a_LC1_A6_aOUT  ;
inv_6091: n_6685  <= TRANSPORT NOT a_N451_aOUT  ;
delay_6092: n_6686  <= TRANSPORT a_N965_aQ  ;
and4_6093: n_6687 <=  n_6688  AND n_6689  AND n_6690  AND n_6691;
delay_6094: n_6688  <= TRANSPORT a_N143_aOUT  ;
delay_6095: n_6689  <= TRANSPORT a_LC1_A6_aOUT  ;
delay_6096: n_6690  <= TRANSPORT a_N451_aOUT  ;
inv_6097: n_6691  <= TRANSPORT NOT a_N965_aQ  ;
and1_6098: n_6692 <=  gnd;
delay_6099: n_6693  <= TRANSPORT nRXC  ;
filter_6100: FILTER_a8251
    PORT MAP (IN1 => n_6693, Y => a_N965_aCLK);
delay_6101: a_N455_aNOT_aOUT  <= TRANSPORT a_N455_aNOT_aIN  ;
xor2_6102: a_N455_aNOT_aIN <=  n_6697  XOR n_6702;
or1_6103: n_6697 <=  n_6698;
and3_6104: n_6698 <=  n_6699  AND n_6700  AND n_6701;
delay_6105: n_6699  <= TRANSPORT a_N390_aOUT  ;
delay_6106: n_6700  <= TRANSPORT a_N451_aOUT  ;
delay_6107: n_6701  <= TRANSPORT a_N965_aQ  ;
and1_6108: n_6702 <=  gnd;
delay_6109: a_N450_aOUT  <= TRANSPORT a_N450_aIN  ;
xor2_6110: a_N450_aIN <=  n_6705  XOR n_6709;
or1_6111: n_6705 <=  n_6706;
and2_6112: n_6706 <=  n_6707  AND n_6708;
delay_6113: n_6707  <= TRANSPORT a_N455_aNOT_aOUT  ;
delay_6114: n_6708  <= TRANSPORT a_N964_aQ  ;
and1_6115: n_6709 <=  gnd;
dff_6116: DFF_a8251
    PORT MAP ( D => a_N963_aD, CLK => a_N963_aCLK, CLRN => a_N963_aCLRN, PRN => vcc,
          Q => a_N963_aQ);
delay_6117: a_N963_aCLRN  <= TRANSPORT nRESET  ;
xor2_6118: a_N963_aD <=  n_6716  XOR n_6727;
or2_6119: n_6716 <=  n_6717  OR n_6722;
and4_6120: n_6717 <=  n_6718  AND n_6719  AND n_6720  AND n_6721;
inv_6121: n_6718  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_6122: n_6719  <= TRANSPORT RXD  ;
inv_6123: n_6720  <= TRANSPORT NOT a_N450_aOUT  ;
delay_6124: n_6721  <= TRANSPORT a_N963_aQ  ;
and4_6125: n_6722 <=  n_6723  AND n_6724  AND n_6725  AND n_6726;
inv_6126: n_6723  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_6127: n_6724  <= TRANSPORT RXD  ;
delay_6128: n_6725  <= TRANSPORT a_N450_aOUT  ;
inv_6129: n_6726  <= TRANSPORT NOT a_N963_aQ  ;
and1_6130: n_6727 <=  gnd;
delay_6131: n_6728  <= TRANSPORT nRXC  ;
filter_6132: FILTER_a8251
    PORT MAP (IN1 => n_6728, Y => a_N963_aCLK);
dff_6133: DFF_a8251
    PORT MAP ( D => a_N964_aD, CLK => a_N964_aCLK, CLRN => a_N964_aCLRN, PRN => vcc,
          Q => a_N964_aQ);
delay_6134: a_N964_aCLRN  <= TRANSPORT nRESET  ;
xor2_6135: a_N964_aD <=  n_6736  XOR n_6747;
or2_6136: n_6736 <=  n_6737  OR n_6742;
and4_6137: n_6737 <=  n_6738  AND n_6739  AND n_6740  AND n_6741;
inv_6138: n_6738  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_6139: n_6739  <= TRANSPORT RXD  ;
delay_6140: n_6740  <= TRANSPORT a_N455_aNOT_aOUT  ;
inv_6141: n_6741  <= TRANSPORT NOT a_N964_aQ  ;
and4_6142: n_6742 <=  n_6743  AND n_6744  AND n_6745  AND n_6746;
inv_6143: n_6743  <= TRANSPORT NOT a_N130_aNOT_aOUT  ;
delay_6144: n_6744  <= TRANSPORT RXD  ;
inv_6145: n_6745  <= TRANSPORT NOT a_N455_aNOT_aOUT  ;
delay_6146: n_6746  <= TRANSPORT a_N964_aQ  ;
and1_6147: n_6747 <=  gnd;
delay_6148: n_6748  <= TRANSPORT nRXC  ;
filter_6149: FILTER_a8251
    PORT MAP (IN1 => n_6748, Y => a_N964_aCLK);
dff_6150: DFF_a8251
    PORT MAP ( D => a_N962_aD, CLK => a_N962_aCLK, CLRN => a_N962_aCLRN, PRN => vcc,
          Q => a_N962_aQ);
delay_6151: a_N962_aCLRN  <= TRANSPORT nRESET  ;
xor2_6152: a_N962_aD <=  n_6756  XOR n_6770;
or3_6153: n_6756 <=  n_6757  OR n_6761  OR n_6765;
and3_6154: n_6757 <=  n_6758  AND n_6759  AND n_6760;
delay_6155: n_6758  <= TRANSPORT a_LC1_A6_aOUT  ;
inv_6156: n_6759  <= TRANSPORT NOT a_N963_aQ  ;
delay_6157: n_6760  <= TRANSPORT a_N962_aQ  ;
and3_6158: n_6761 <=  n_6762  AND n_6763  AND n_6764;
delay_6159: n_6762  <= TRANSPORT a_LC1_A6_aOUT  ;
inv_6160: n_6763  <= TRANSPORT NOT a_N450_aOUT  ;
delay_6161: n_6764  <= TRANSPORT a_N962_aQ  ;
and4_6162: n_6765 <=  n_6766  AND n_6767  AND n_6768  AND n_6769;
delay_6163: n_6766  <= TRANSPORT a_LC1_A6_aOUT  ;
delay_6164: n_6767  <= TRANSPORT a_N450_aOUT  ;
delay_6165: n_6768  <= TRANSPORT a_N963_aQ  ;
inv_6166: n_6769  <= TRANSPORT NOT a_N962_aQ  ;
and1_6167: n_6770 <=  gnd;
delay_6168: n_6771  <= TRANSPORT nRXC  ;
filter_6169: FILTER_a8251
    PORT MAP (IN1 => n_6771, Y => a_N962_aCLK);
delay_6170: a_LC7_C15_aOUT  <= TRANSPORT a_LC7_C15_aIN  ;
xor2_6171: a_LC7_C15_aIN <=  n_6775  XOR n_6783;
or2_6172: n_6775 <=  n_6776  OR n_6780;
and3_6173: n_6776 <=  n_6777  AND n_6778  AND n_6779;
inv_6174: n_6777  <= TRANSPORT NOT a_N1120_aNOT_aOUT  ;
inv_6175: n_6778  <= TRANSPORT NOT a_N1121_aNOT_aOUT  ;
delay_6176: n_6779  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and2_6177: n_6780 <=  n_6781  AND n_6782;
delay_6178: n_6781  <= TRANSPORT a_N613_aOUT  ;
delay_6179: n_6782  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_6180: n_6783 <=  gnd;
dff_6181: DFF_a8251
    PORT MAP ( D => a_SCMND_OUT_F2_G_aD, CLK => a_SCMND_OUT_F2_G_aCLK, CLRN => a_SCMND_OUT_F2_G_aCLRN,
          PRN => vcc, Q => a_SCMND_OUT_F2_G_aQ);
delay_6182: a_SCMND_OUT_F2_G_aCLRN  <= TRANSPORT nRESET  ;
xor2_6183: a_SCMND_OUT_F2_G_aD <=  n_6790  XOR n_6798;
or2_6184: n_6790 <=  n_6791  OR n_6794;
and2_6185: n_6791 <=  n_6792  AND n_6793;
delay_6186: n_6792  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_6187: n_6793  <= TRANSPORT a_LC7_C15_aOUT  ;
and3_6188: n_6794 <=  n_6795  AND n_6796  AND n_6797;
delay_6189: n_6795  <= TRANSPORT a_N82_aNOT_aOUT  ;
delay_6190: n_6796  <= TRANSPORT DIN(2)  ;
delay_6191: n_6797  <= TRANSPORT a_N701_aNOT_aOUT  ;
and1_6192: n_6798 <=  gnd;
delay_6193: n_6799  <= TRANSPORT CLK  ;
filter_6194: FILTER_a8251
    PORT MAP (IN1 => n_6799, Y => a_SCMND_OUT_F2_G_aCLK);
delay_6195: a_N659_aNOT_aOUT  <= TRANSPORT a_N659_aNOT_aIN  ;
xor2_6196: a_N659_aNOT_aIN <=  n_6803  XOR n_6808;
or1_6197: n_6803 <=  n_6804;
and3_6198: n_6804 <=  n_6805  AND n_6806  AND n_6807;
inv_6199: n_6805  <= TRANSPORT NOT a_N735_aNOT_aOUT  ;
inv_6200: n_6806  <= TRANSPORT NOT RXD  ;
delay_6201: n_6807  <= TRANSPORT a_SCMND_OUT_F2_G_aQ  ;
and1_6202: n_6808 <=  gnd;
delay_6203: a_LC4_D12_aOUT  <= TRANSPORT a_LC4_D12_aIN  ;
xor2_6204: a_LC4_D12_aIN <=  n_6811  XOR n_6818;
or2_6205: n_6811 <=  n_6812  OR n_6815;
and2_6206: n_6812 <=  n_6813  AND n_6814;
inv_6207: n_6813  <= TRANSPORT NOT a_N1152_aNOT_aOUT  ;
inv_6208: n_6814  <= TRANSPORT NOT a_N63_aQ  ;
and2_6209: n_6815 <=  n_6816  AND n_6817;
inv_6210: n_6816  <= TRANSPORT NOT a_N1152_aNOT_aOUT  ;
inv_6211: n_6817  <= TRANSPORT NOT a_N62_aQ  ;
and1_6212: n_6818 <=  gnd;
delay_6213: a_LC8_D12_aOUT  <= TRANSPORT a_LC8_D12_aIN  ;
xor2_6214: a_LC8_D12_aIN <=  n_6821  XOR n_6827;
or1_6215: n_6821 <=  n_6822;
and4_6216: n_6822 <=  n_6823  AND n_6824  AND n_6825  AND n_6826;
inv_6217: n_6823  <= TRANSPORT NOT a_N1183_aNOT_aOUT  ;
delay_6218: n_6824  <= TRANSPORT a_N1164_aOUT  ;
delay_6219: n_6825  <= TRANSPORT a_N62_aQ  ;
inv_6220: n_6826  <= TRANSPORT NOT a_N63_aQ  ;
and1_6221: n_6827 <=  gnd;
delay_6222: a_LC6_D12_aOUT  <= TRANSPORT a_LC6_D12_aIN  ;
xor2_6223: a_LC6_D12_aIN <=  n_6830  XOR n_6838;
or3_6224: n_6830 <=  n_6831  OR n_6834  OR n_6836;
and2_6225: n_6831 <=  n_6832  AND n_6833;
delay_6226: n_6832  <= TRANSPORT a_N1158_aOUT  ;
delay_6227: n_6833  <= TRANSPORT a_N659_aNOT_aOUT  ;
and1_6228: n_6834 <=  n_6835;
delay_6229: n_6835  <= TRANSPORT a_LC4_D12_aOUT  ;
and1_6230: n_6836 <=  n_6837;
delay_6231: n_6837  <= TRANSPORT a_LC8_D12_aOUT  ;
and1_6232: n_6838 <=  gnd;
delay_6233: a_LC7_D12_aOUT  <= TRANSPORT a_LC7_D12_aIN  ;
xor2_6234: a_LC7_D12_aIN <=  n_6841  XOR n_6849;
or3_6235: n_6841 <=  n_6842  OR n_6845  OR n_6847;
and2_6236: n_6842 <=  n_6843  AND n_6844;
inv_6237: n_6843  <= TRANSPORT NOT a_N132_aOUT  ;
delay_6238: n_6844  <= TRANSPORT a_N1080_aOUT  ;
and1_6239: n_6845 <=  n_6846;
delay_6240: n_6846  <= TRANSPORT a_LC6_D12_aOUT  ;
and1_6241: n_6847 <=  n_6848;
inv_6242: n_6848  <= TRANSPORT NOT a_N155_aOUT  ;
and1_6243: n_6849 <=  gnd;
dff_6244: DFF_a8251
    PORT MAP ( D => a_N61_aD, CLK => a_N61_aCLK, CLRN => a_N61_aCLRN, PRN => vcc,
          Q => a_N61_aQ);
delay_6245: a_N61_aCLRN  <= TRANSPORT nRESET  ;
xor2_6246: a_N61_aD <=  n_6856  XOR n_6866;
or3_6247: n_6856 <=  n_6857  OR n_6860  OR n_6863;
and2_6248: n_6857 <=  n_6858  AND n_6859;
inv_6249: n_6858  <= TRANSPORT NOT a_N83_aOUT  ;
delay_6250: n_6859  <= TRANSPORT a_N1067_aOUT  ;
and2_6251: n_6860 <=  n_6861  AND n_6862;
inv_6252: n_6861  <= TRANSPORT NOT a_N83_aOUT  ;
delay_6253: n_6862  <= TRANSPORT a_N91_aOUT  ;
and2_6254: n_6863 <=  n_6864  AND n_6865;
inv_6255: n_6864  <= TRANSPORT NOT a_N83_aOUT  ;
delay_6256: n_6865  <= TRANSPORT a_LC7_D12_aOUT  ;
and1_6257: n_6866 <=  gnd;
delay_6258: n_6867  <= TRANSPORT nRXC  ;
filter_6259: FILTER_a8251
    PORT MAP (IN1 => n_6867, Y => a_N61_aCLK);
delay_6260: a_LC2_D11_aOUT  <= TRANSPORT a_LC2_D11_aIN  ;
xor2_6261: a_LC2_D11_aIN <=  n_6871  XOR n_6876;
or1_6262: n_6871 <=  n_6872;
and3_6263: n_6872 <=  n_6873  AND n_6874  AND n_6875;
inv_6264: n_6873  <= TRANSPORT NOT a_LC2_D19_aOUT  ;
delay_6265: n_6874  <= TRANSPORT a_N64_aQ  ;
inv_6266: n_6875  <= TRANSPORT NOT a_N61_aQ  ;
and1_6267: n_6876 <=  gnd;
delay_6268: a_N653_aOUT  <= TRANSPORT a_N653_aIN  ;
xor2_6269: a_N653_aIN <=  n_6879  XOR n_6887;
or2_6270: n_6879 <=  n_6880  OR n_6884;
and3_6271: n_6880 <=  n_6881  AND n_6882  AND n_6883;
delay_6272: n_6881  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_6273: n_6882  <= TRANSPORT a_N134_aNOT_aOUT  ;
delay_6274: n_6883  <= TRANSPORT a_LC6_A13_aOUT  ;
and2_6275: n_6884 <=  n_6885  AND n_6886;
delay_6276: n_6885  <= TRANSPORT a_LC6_A13_aOUT  ;
inv_6277: n_6886  <= TRANSPORT NOT a_N1555_aQ  ;
and1_6278: n_6887 <=  gnd;
delay_6279: a_N655_aOUT  <= TRANSPORT a_N655_aIN  ;
xor2_6280: a_N655_aIN <=  n_6889  XOR n_6897;
or3_6281: n_6889 <=  n_6890  OR n_6892  OR n_6895;
and1_6282: n_6890 <=  n_6891;
delay_6283: n_6891  <= TRANSPORT a_N653_aOUT  ;
and2_6284: n_6892 <=  n_6893  AND n_6894;
delay_6285: n_6893  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_6286: n_6894  <= TRANSPORT a_N1193_aOUT  ;
and1_6287: n_6895 <=  n_6896;
inv_6288: n_6896  <= TRANSPORT NOT a_N1037_aNOT_aOUT  ;
and1_6289: n_6897 <=  gnd;
delay_6290: a_N75_aOUT  <= TRANSPORT a_N75_aIN  ;
xor2_6291: a_N75_aIN <=  n_6900  XOR n_6907;
or2_6292: n_6900 <=  n_6901  OR n_6904;
and2_6293: n_6901 <=  n_6902  AND n_6903;
delay_6294: n_6902  <= TRANSPORT EXTSYNCD  ;
delay_6295: n_6903  <= TRANSPORT a_SMODE_OUT_F6_G_aQ  ;
and2_6296: n_6904 <=  n_6905  AND n_6906;
delay_6297: n_6905  <= TRANSPORT a_N655_aOUT  ;
inv_6298: n_6906  <= TRANSPORT NOT a_SMODE_OUT_F6_G_aQ  ;
and1_6299: n_6907 <=  gnd;
delay_6300: a_LC3_D18_aOUT  <= TRANSPORT a_LC3_D18_aIN  ;
xor2_6301: a_LC3_D18_aIN <=  n_6910  XOR n_6916;
or1_6302: n_6910 <=  n_6911;
and4_6303: n_6911 <=  n_6912  AND n_6913  AND n_6914  AND n_6915;
inv_6304: n_6912  <= TRANSPORT NOT a_N1118_aNOT_aOUT  ;
delay_6305: n_6913  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_6306: n_6914  <= TRANSPORT a_N64_aQ  ;
inv_6307: n_6915  <= TRANSPORT NOT a_N62_aQ  ;
and1_6308: n_6916 <=  gnd;
delay_6309: a_LC2_D8_aOUT  <= TRANSPORT a_LC2_D8_aIN  ;
xor2_6310: a_LC2_D8_aIN <=  n_6919  XOR n_6932;
or4_6311: n_6919 <=  n_6920  OR n_6923  OR n_6926  OR n_6929;
and2_6312: n_6920 <=  n_6921  AND n_6922;
delay_6313: n_6921  <= TRANSPORT a_LC3_D18_aOUT  ;
inv_6314: n_6922  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_6315: n_6923 <=  n_6924  AND n_6925;
delay_6316: n_6924  <= TRANSPORT a_N132_aOUT  ;
delay_6317: n_6925  <= TRANSPORT a_LC3_D18_aOUT  ;
and2_6318: n_6926 <=  n_6927  AND n_6928;
delay_6319: n_6927  <= TRANSPORT a_N1080_aOUT  ;
inv_6320: n_6928  <= TRANSPORT NOT a_SMODE_OUT_F4_G_aQ  ;
and2_6321: n_6929 <=  n_6930  AND n_6931;
delay_6322: n_6930  <= TRANSPORT a_N132_aOUT  ;
delay_6323: n_6931  <= TRANSPORT a_N1080_aOUT  ;
and1_6324: n_6932 <=  gnd;
delay_6325: a_LC7_D8_aNOT_aOUT  <= TRANSPORT a_LC7_D8_aNOT_aIN  ;
xor2_6326: a_LC7_D8_aNOT_aIN <=  n_6935  XOR n_6939;
or1_6327: n_6935 <=  n_6936;
and2_6328: n_6936 <=  n_6937  AND n_6938;
inv_6329: n_6937  <= TRANSPORT NOT a_N1149_aNOT_aOUT  ;
inv_6330: n_6938  <= TRANSPORT NOT a_N64_aQ  ;
and1_6331: n_6939 <=  gnd;
delay_6332: a_N656_aNOT_aOUT  <= TRANSPORT a_N656_aNOT_aIN  ;
xor2_6333: a_N656_aNOT_aIN <=  n_6942  XOR n_6951;
or2_6334: n_6942 <=  n_6943  OR n_6947;
and3_6335: n_6943 <=  n_6944  AND n_6945  AND n_6946;
inv_6336: n_6944  <= TRANSPORT NOT RXD  ;
delay_6337: n_6945  <= TRANSPORT a_LC7_D8_aNOT_aOUT  ;
delay_6338: n_6946  <= TRANSPORT a_N63_aQ  ;
and3_6339: n_6947 <=  n_6948  AND n_6949  AND n_6950;
delay_6340: n_6948  <= TRANSPORT a_N1120_aNOT_aOUT  ;
delay_6341: n_6949  <= TRANSPORT a_LC7_D8_aNOT_aOUT  ;
inv_6342: n_6950  <= TRANSPORT NOT a_N63_aQ  ;
and1_6343: n_6951 <=  gnd;
delay_6344: a_LC5_D8_aOUT  <= TRANSPORT a_LC5_D8_aIN  ;
xor2_6345: a_LC5_D8_aIN <=  n_6954  XOR n_6963;
or4_6346: n_6954 <=  n_6955  OR n_6957  OR n_6959  OR n_6961;
and1_6347: n_6955 <=  n_6956;
delay_6348: n_6956  <= TRANSPORT a_LC2_D8_aOUT  ;
and1_6349: n_6957 <=  n_6958;
delay_6350: n_6958  <= TRANSPORT a_N656_aNOT_aOUT  ;
and1_6351: n_6959 <=  n_6960;
delay_6352: n_6960  <= TRANSPORT a_N1069_aOUT  ;
and1_6353: n_6961 <=  n_6962;
inv_6354: n_6962  <= TRANSPORT NOT a_N125_aOUT  ;
and1_6355: n_6963 <=  gnd;
delay_6356: a_LC3_D12_aOUT  <= TRANSPORT a_LC3_D12_aIN  ;
xor2_6357: a_LC3_D12_aIN <=  n_6966  XOR n_6975;
or4_6358: n_6966 <=  n_6967  OR n_6969  OR n_6971  OR n_6973;
and1_6359: n_6967 <=  n_6968;
delay_6360: n_6968  <= TRANSPORT a_LC5_D8_aOUT  ;
and1_6361: n_6969 <=  n_6970;
delay_6362: n_6970  <= TRANSPORT a_N1067_aOUT  ;
and1_6363: n_6971 <=  n_6972;
delay_6364: n_6972  <= TRANSPORT a_N91_aOUT  ;
and1_6365: n_6973 <=  n_6974;
delay_6366: n_6974  <= TRANSPORT a_N659_aNOT_aOUT  ;
and1_6367: n_6975 <=  gnd;
delay_6368: a_LC5_D12_aOUT  <= TRANSPORT a_LC5_D12_aIN  ;
xor2_6369: a_LC5_D12_aIN <=  n_6978  XOR n_6986;
or3_6370: n_6978 <=  n_6979  OR n_6981  OR n_6984;
and1_6371: n_6979 <=  n_6980;
delay_6372: n_6980  <= TRANSPORT a_LC3_D12_aOUT  ;
and2_6373: n_6981 <=  n_6982  AND n_6983;
delay_6374: n_6982  <= TRANSPORT a_N95_aNOT_aOUT  ;
delay_6375: n_6983  <= TRANSPORT a_LC7_D7_aOUT  ;
and1_6376: n_6984 <=  n_6985;
delay_6377: n_6985  <= TRANSPORT a_N108_aNOT_aOUT  ;
and1_6378: n_6986 <=  gnd;
dff_6379: DFF_a8251
    PORT MAP ( D => a_N63_aD, CLK => a_N63_aCLK, CLRN => a_N63_aCLRN, PRN => vcc,
          Q => a_N63_aQ);
delay_6380: a_N63_aCLRN  <= TRANSPORT nRESET  ;
xor2_6381: a_N63_aD <=  n_6993  XOR n_7001;
or2_6382: n_6993 <=  n_6994  OR n_6998;
and3_6383: n_6994 <=  n_6995  AND n_6996  AND n_6997;
inv_6384: n_6995  <= TRANSPORT NOT a_N83_aOUT  ;
delay_6385: n_6996  <= TRANSPORT a_LC2_D11_aOUT  ;
delay_6386: n_6997  <= TRANSPORT a_N75_aOUT  ;
and2_6387: n_6998 <=  n_6999  AND n_7000;
inv_6388: n_6999  <= TRANSPORT NOT a_N83_aOUT  ;
delay_6389: n_7000  <= TRANSPORT a_LC5_D12_aOUT  ;
and1_6390: n_7001 <=  gnd;
delay_6391: n_7002  <= TRANSPORT nRXC  ;
filter_6392: FILTER_a8251
    PORT MAP (IN1 => n_7002, Y => a_N63_aCLK);
delay_6393: a_LC1_C2_aOUT  <= TRANSPORT a_LC1_C2_aIN  ;
xor2_6394: a_LC1_C2_aIN <=  n_7005  XOR n_7011;
or1_6395: n_7005 <=  n_7006;
and4_6396: n_7006 <=  n_7007  AND n_7008  AND n_7009  AND n_7010;
delay_6397: n_7007  <= TRANSPORT a_N82_aNOT_aOUT  ;
inv_6398: n_7008  <= TRANSPORT NOT a_N1754_aQ  ;
inv_6399: n_7009  <= TRANSPORT NOT a_N1757_aQ  ;
inv_6400: n_7010  <= TRANSPORT NOT a_N1756_aQ  ;
and1_6401: n_7011 <=  gnd;

END REVISION1_2;
